//: version "1.8.7"

module CLL(G3, P1, G1, G0, Cin, G2, P2, PG, C2, C4, C1, P3, P0, GG, C3);
//: interface  /sz:(974, 86) /bd:[ Ti0>P3(120/974) Ti1>G3(182/974) Ti2>P2(402/974) Ti3>G2(457/974) Ti4>P1(657/974) Ti5>G1(710/974) Ti6>P0(887/974) Ti7>G0(946/974) Ri0>Cin(57/86) To0<C3(242/974) To1<C2(505/974) To2<C1(746/974) Lo0<C4(45/86) Bo0<PG(685/974) Bo1<GG(837/974) ]
input G2;    //: /sn:0 {0}(297,703)(267,703){1}
//: {2}(265,701)(265,518){3}
//: {4}(267,516)(362,516){5}
//: {6}(263,516)(167,516){7}
//: {8}(265,705)(265,851)(299,851){9}
output GG;    //: /sn:0 {0}(427,807)(398,807){1}
input P1;    //: /sn:0 {0}(300,782)(243,782)(243,742){1}
//: {2}(245,740)(299,740){3}
//: {4}(243,738)(243,634){5}
//: {6}(245,632)(298,632){7}
//: {8}(243,630)(243,590){9}
//: {10}(245,588)(298,588){11}
//: {12}(243,586)(243,523)(216,523)(216,506){13}
//: {14}(218,504)(286,504){15}
//: {16}(216,502)(216,474){17}
//: {18}(218,472)(287,472){19}
//: {20}(216,470)(216,410){21}
//: {22}(218,408)(286,408){23}
//: {24}(216,406)(216,374){25}
//: {26}(218,372)(287,372){27}
//: {28}(214,372)(166,372){29}
output C3;    //: /sn:0 {0}(408,508)(383,508){1}
output PG;    //: /sn:0 /dp:1 {0}(320,742)(364,742){1}
input G0;    //: /sn:0 /dp:1 {0}(334,261)(261,261)(261,294)(211,294){1}
//: {2}(207,294)(177,294)(177,309)(167,309){3}
//: {4}(209,296)(209,411){5}
//: {6}(211,413)(286,413){7}
//: {8}(209,415)(209,497){9}
//: {10}(211,499)(286,499){11}
//: {12}(209,501)(209,625){13}
//: {14}(211,627)(298,627){15}
//: {16}(209,629)(209,777)(300,777){17}
output C4;    //: /sn:0 {0}(438,655)(403,655){1}
output C2;    //: /sn:0 {0}(401,385)(369,385){1}
input Cin;    //: /sn:0 /dp:7 {0}(287,362)(232,362){1}
//: {2}(230,360)(230,287){3}
//: {4}(230,283)(230,258)(235,258){5}
//: {6}(228,285)(167,285){7}
//: {8}(230,364)(230,460){9}
//: {10}(232,462)(287,462){11}
//: {12}(230,464)(230,578)(298,578){13}
input P3;    //: /sn:0 /dp:1 {0}(299,745)(260,745){1}
//: {2}(258,743)(258,710){3}
//: {4}(260,708)(297,708){5}
//: {6}(258,706)(258,680){7}
//: {8}(260,678)(298,678){9}
//: {10}(258,676)(258,644){11}
//: {12}(260,642)(298,642){13}
//: {14}(258,640)(258,600){15}
//: {16}(260,598)(298,598){17}
//: {18}(256,598)(170,598)(170,598)(167,598){19}
//: {20}(258,747)(258,790){21}
//: {22}(260,792)(300,792){23}
//: {24}(258,794)(258,824){25}
//: {26}(260,826)(300,826){27}
//: {28}(258,828)(258,856)(299,856){29}
input G1;    //: /sn:0 {0}(166,385)(200,385){1}
//: {2}(204,385)(348,385){3}
//: {4}(202,387)(202,511){5}
//: {6}(204,513)(279,513)(279,536)(289,536){7}
//: {8}(202,515)(202,666){9}
//: {10}(204,668)(298,668){11}
//: {12}(202,670)(202,816)(300,816){13}
input G3;    //: /sn:0 /dp:1 {0}(382,655)(224,655){1}
//: {2}(220,655)(166,655){3}
//: {4}(222,657)(222,805)(377,805){5}
output C1;    //: /sn:0 /dp:1 {0}(355,259)(399,259){1}
input P0;    //: /sn:0 {0}(287,467)(238,467){1}
//: {2}(236,465)(236,369){3}
//: {4}(238,367)(287,367){5}
//: {6}(234,367)(221,367)(221,236){7}
//: {8}(223,234)(229,234)(229,253)(235,253){9}
//: {10}(219,234)(180,234)(180,234)(166,234){11}
//: {12}(236,469)(236,581){13}
//: {14}(238,583)(298,583){15}
//: {16}(236,585)(236,735)(299,735){17}
input P2;    //: /sn:0 {0}(299,750)(275,750){1}
//: {2}(273,748)(273,675){3}
//: {4}(275,673)(298,673){5}
//: {6}(271,673)(250,673)(250,639){7}
//: {8}(252,637)(298,637){9}
//: {10}(250,635)(250,595){11}
//: {12}(252,593)(298,593){13}
//: {14}(250,591)(250,511){15}
//: {16}(252,509)(286,509){17}
//: {18}(248,509)(227,509){19}
//: {20}(225,507)(225,479){21}
//: {22}(227,477)(287,477){23}
//: {24}(223,477)(168,477){25}
//: {26}(225,511)(225,541)(289,541){27}
//: {28}(273,752)(273,785){29}
//: {30}(275,787)(300,787){31}
//: {32}(273,789)(273,821)(300,821){33}
wire w6;    //: /sn:0 {0}(320,854)(367,854)(367,815)(377,815){1}
wire w4;    //: /sn:0 {0}(321,784)(367,784)(367,800)(377,800){1}
wire w39;    //: /sn:0 /dp:1 {0}(318,706)(345,706)(345,665)(382,665){1}
wire w3;    //: /sn:0 {0}(307,411)(338,411)(338,390)(348,390){1}
wire D8;    //: /sn:0 {0}(308,367)(338,367)(338,380)(348,380){1}
wire w42;    //: /sn:0 /dp:1 {0}(319,588)(346,588)(346,645)(382,645){1}
wire w18;    //: /sn:0 /dp:1 {0}(307,504)(317,504)(317,506)(362,506){1}
wire w8;    //: /sn:0 {0}(377,810)(359,810)(359,821)(321,821){1}
wire w44;    //: /sn:0 {0}(362,511)(320,511)(320,539)(310,539){1}
wire w45;    //: /sn:0 /dp:1 {0}(308,469)(321,469)(321,501)(362,501){1}
wire w2;    //: /sn:0 /dp:1 {0}(256,256)(334,256){1}
wire w15;    //: /sn:0 /dp:1 {0}(319,634)(340,634)(340,650)(382,650){1}
wire w40;    //: /sn:0 /dp:1 {0}(319,673)(339,673)(339,660)(382,660){1}
//: enddecls

  and g44 (.I0(G1), .I1(P2), .I2(P3), .Z(w40));   //: @(309,673) /sn:0 /delay:" 3" /w:[ 11 5 9 0 ]
  //: input g8 (G3) @(164,655) /sn:0 /w:[ 3 ]
  //: input g4 (P1) @(164,372) /sn:0 /w:[ 29 ]
  //: joint g47 (P3) @(258, 642) /w:[ 12 14 -1 11 ]
  //: joint g16 (Cin) @(230, 285) /w:[ -1 4 6 3 ]
  //: input g3 (G1) @(164,385) /sn:0 /w:[ 0 ]
  //: joint g17 (P0) @(221, 234) /w:[ 8 -1 10 7 ]
  and g26 (.I0(G0), .I1(P1), .I2(P2), .Z(w18));   //: @(297,504) /sn:0 /delay:" 3" /w:[ 11 15 17 0 ]
  //: input g2 (G0) @(165,309) /sn:0 /w:[ 3 ]
  //: joint g23 (Cin) @(230, 362) /w:[ 1 2 -1 8 ]
  and g30 (.I0(G1), .I1(P2), .Z(w44));   //: @(300,539) /sn:0 /delay:" 3" /w:[ 7 27 1 ]
  //: joint g24 (P0) @(236, 367) /w:[ 4 -1 6 3 ]
  and g39 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w15));   //: @(309,634) /sn:0 /delay:" 3" /w:[ 15 7 9 13 0 ]
  //: input g1 (Cin) @(165,285) /sn:0 /w:[ 7 ]
  //: joint g60 (G0) @(209, 627) /w:[ 14 13 -1 16 ]
  //: joint g29 (P2) @(225, 477) /w:[ 22 -1 24 21 ]
  or g51 (.I0(w42), .I1(w15), .I2(G3), .I3(w40), .I4(w39), .Z(C4));   //: @(393,655) /sn:0 /delay:" 3" /w:[ 1 1 0 1 1 1 ]
  //: joint g70 (P3) @(258, 826) /w:[ 26 25 -1 28 ]
  and g18 (.I0(P1), .I1(G0), .Z(w3));   //: @(297,411) /sn:0 /delay:" 3" /w:[ 23 7 0 ]
  //: joint g65 (G1) @(202, 668) /w:[ 10 9 -1 12 ]
  //: joint g25 (P1) @(216, 408) /w:[ 22 24 -1 21 ]
  or g10 (.I0(w2), .I1(G0), .Z(C1));   //: @(345,259) /sn:0 /delay:" 3" /w:[ 1 0 0 ]
  and g64 (.I0(G1), .I1(P2), .I2(P3), .Z(w8));   //: @(311,821) /sn:0 /delay:" 3" /w:[ 13 33 27 1 ]
  //: joint g72 (G3) @(222, 655) /w:[ 1 -1 2 4 ]
  //: joint g49 (G2) @(265, 516) /w:[ 4 -1 6 3 ]
  //: joint g50 (P3) @(258, 678) /w:[ 8 10 -1 7 ]
  //: input g6 (G2) @(165,516) /sn:0 /w:[ 7 ]
  and g68 (.I0(G2), .I1(P3), .Z(w6));   //: @(310,854) /sn:0 /delay:" 3" /w:[ 9 29 0 ]
  //: joint g58 (P3) @(258, 708) /w:[ 4 6 -1 3 ]
  //: joint g56 (P1) @(243, 632) /w:[ 6 8 -1 5 ]
  //: joint g35 (Cin) @(230, 462) /w:[ 10 9 -1 12 ]
  and g9 (.I0(P0), .I1(Cin), .Z(w2));   //: @(246,256) /sn:0 /delay:" 3" /w:[ 9 5 0 ]
  //: input g7 (P2) @(166,477) /sn:0 /w:[ 25 ]
  and g73 (.I0(P0), .I1(P1), .I2(P3), .I3(P2), .Z(PG));   //: @(310,742) /sn:0 /delay:" 3" /w:[ 17 3 0 0 0 ]
  or g71 (.I0(w4), .I1(G3), .I2(w8), .I3(w6), .Z(GG));   //: @(388,807) /sn:0 /delay:" 3" /w:[ 1 5 0 1 1 ]
  and g59 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w4));   //: @(311,784) /sn:0 /delay:" 3" /w:[ 17 0 31 23 0 ]
  //: joint g31 (G1) @(202, 385) /w:[ 2 -1 1 4 ]
  and g22 (.I0(Cin), .I1(P0), .I2(P1), .I3(P2), .Z(w45));   //: @(298,469) /sn:0 /delay:" 3" /w:[ 11 0 19 23 0 ]
  //: joint g67 (P3) @(258, 792) /w:[ 22 21 -1 24 ]
  //: joint g45 (G1) @(202, 513) /w:[ 6 5 -1 8 ]
  //: joint g41 (P1) @(243, 588) /w:[ 10 12 -1 9 ]
  //: joint g36 (P0) @(236, 467) /w:[ 1 2 -1 12 ]
  or g33 (.I0(w45), .I1(w18), .I2(w44), .I3(G2), .Z(C3));   //: @(373,508) /sn:0 /delay:" 3" /w:[ 1 1 0 5 1 ]
  //: joint g54 (P0) @(236, 583) /w:[ 14 13 -1 16 ]
  //: joint g69 (G2) @(265, 703) /w:[ 1 2 -1 8 ]
  //: output g52 (PG) @(361,742) /sn:0 /w:[ 1 ]
  //: joint g42 (P2) @(250, 593) /w:[ 12 14 -1 11 ]
  //: joint g40 (G0) @(209, 499) /w:[ 10 9 -1 12 ]
  //: joint g66 (P2) @(273, 787) /w:[ 30 29 -1 32 ]
  //: output g12 (C2) @(398,385) /sn:0 /w:[ 0 ]
  //: joint g57 (P2) @(273, 673) /w:[ 4 -1 6 3 ]
  //: joint g46 (P2) @(250, 637) /w:[ 8 10 -1 7 ]
  //: joint g28 (P1) @(216, 472) /w:[ 18 20 -1 17 ]
  and g34 (.I0(Cin), .I1(P0), .I2(P1), .I3(P2), .I4(P3), .Z(w42));   //: @(309,588) /sn:0 /anc:1 /delay:" 3" /w:[ 13 15 11 13 17 0 ]
  //: output g14 (C4) @(435,655) /sn:0 /w:[ 0 ]
  //: output g11 (C1) @(396,259) /sn:0 /w:[ 1 ]
  //: input g5 (P3) @(165,598) /sn:0 /w:[ 19 ]
  //: joint g19 (P1) @(216, 372) /w:[ 26 -1 28 25 ]
  or g21 (.I0(D8), .I1(G1), .I2(w3), .Z(C2));   //: @(359,385) /sn:0 /delay:" 3" /w:[ 1 3 1 1 ]
  //: joint g61 (P3) @(258, 745) /w:[ 1 2 -1 20 ]
  //: joint g32 (P1) @(216, 504) /w:[ 14 16 -1 13 ]
  //: joint g20 (G0) @(209, 294) /w:[ 1 -1 2 4 ]
  //: joint g43 (P3) @(258, 598) /w:[ 16 -1 18 15 ]
  //: joint g38 (P2) @(250, 509) /w:[ 16 -1 18 15 ]
  and g15 (.I0(Cin), .I1(P0), .I2(P1), .Z(D8));   //: @(298,367) /sn:0 /delay:" 3" /w:[ 0 5 27 0 ]
  //: input g0 (P0) @(164,234) /sn:0 /w:[ 11 ]
  //: joint g27 (G0) @(209, 413) /w:[ 6 5 -1 8 ]
  and g48 (.I0(G2), .I1(P3), .Z(w39));   //: @(308,706) /sn:0 /delay:" 3" /w:[ 0 5 0 ]
  //: joint g37 (P2) @(225, 509) /w:[ 19 20 -1 26 ]
  //: joint g62 (P2) @(273, 750) /w:[ 1 2 -1 28 ]
  //: joint g55 (P1) @(243, 740) /w:[ 2 4 -1 1 ]
  //: output g53 (GG) @(424,807) /sn:0 /w:[ 0 ]
  //: output g13 (C3) @(405,508) /sn:0 /w:[ 0 ]

endmodule

module CLA16Bits(B, Cin, A, GG, Cout, PG, S);
//: interface  /sz:(322, 143) /bd:[ Ti0>A[15:0](70/322) Ti1>B[15:0](209/322) Ri0>Cin(75/143) Lo0<PG(111/143) Lo1<GG(58/143) Bo0<Cout(182/322) Bo1<S[15:0](235/322) ]
input [15:0] B;    //: /sn:0 {0}(-203,-33)(-70,-33){1}
//: {2}(-69,-33)(191,-33){3}
//: {4}(192,-33)(463,-33){5}
//: {6}(464,-33)(723,-33){7}
//: {8}(724,-33)(877,-33){9}
output GG;    //: /sn:0 /dp:1 {0}(693,354)(693,421){1}
input [15:0] A;    //: /sn:0 {0}(875,-108)(686,-108){1}
//: {2}(685,-108)(415,-108){3}
//: {4}(414,-108)(157,-108){5}
//: {6}(156,-108)(-107,-108){7}
//: {8}(-108,-108)(-201,-108){9}
output PG;    //: /sn:0 /dp:1 {0}(541,354)(541,419){1}
input Cin;    //: /sn:0 {0}(826,93)(971,93)(971,94){1}
//: {2}(973,96)(979,96)(979,87)(989,87){3}
//: {4}(971,98)(971,324)(831,324){5}
output Cout;    //: /sn:0 /dp:1 {0}(-145,312)(-265,312)(-265,316)(-255,316){1}
output [15:0] S;    //: /sn:0 /dp:1 {0}(885,194)(925,194){1}
wire w16;    //: /sn:0 {0}(802,266)(802,232)(750,232)(750,156){1}
wire w6;    //: /sn:0 {0}(294,90)(361,90)(361,266){1}
wire [3:0] w7;    //: /sn:0 {0}(155,153)(155,189)(879,189){1}
wire w25;    //: /sn:0 /dp:1 {0}(98,266)(98,82)(32,82){1}
wire [3:0] w39;    //: /sn:0 {0}(687,156)(687,209)(879,209){1}
wire w22;    //: /sn:0 {0}(38,266)(38,223)(-44,223)(-44,145){1}
wire [3:0] w0;    //: /sn:0 /dp:1 {0}(157,-104)(157,-83)(155,-83)(155,55){1}
wire [3:0] w36;    //: /sn:0 {0}(687,58)(687,46)(686,46)(686,-104){1}
wire w20;    //: /sn:0 {0}(313,266)(313,234)(218,234)(218,153){1}
wire [3:0] w37;    //: /sn:0 {0}(724,58)(724,-29){1}
wire w18;    //: /sn:0 {0}(566,266)(566,252)(486,252)(486,157){1}
wire w19;    //: /sn:0 {0}(513,266)(513,167)(529,167)(529,157){1}
wire w12;    //: /sn:0 {0}(562,94)(602,94)(602,266){1}
wire w23;    //: /sn:0 {0}(-24,266)(-24,250)(-1,250)(-1,145){1}
wire [3:0] w10;    //: /sn:0 {0}(423,59)(423,33)(415,33)(415,-104){1}
wire [3:0] w1;    //: /sn:0 /dp:1 {0}(192,-29)(192,55){1}
wire [3:0] w31;    //: /sn:0 /dp:1 {0}(879,199)(423,199)(423,157){1}
wire w17;    //: /sn:0 {0}(743,266)(743,241)(791,241)(791,156){1}
wire [3:0] w27;    //: /sn:0 /dp:1 {0}(464,-29)(464,49)(460,49)(460,59){1}
wire [3:0] w14;    //: /sn:0 /dp:1 {0}(-107,-104)(-107,47){1}
wire [3:0] w2;    //: /sn:0 {0}(-70,47)(-70,-21)(-69,-21)(-69,-29){1}
wire [3:0] w26;    //: /sn:0 /dp:1 {0}(879,179)(-107,179)(-107,145){1}
wire w9;    //: /sn:0 /dp:1 {0}(261,153)(261,256)(258,256)(258,266){1}
//: enddecls

  CLL g4 (.P3(w23), .G3(w22), .P2(w9), .G2(w20), .P1(w19), .G1(w18), .P0(w17), .G0(w16), .Cin(Cin), .C3(w25), .C2(w6), .C1(w12), .C4(Cout), .PG(PG), .GG(GG));   //: @(-144, 267) /sz:(974, 86) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>5 To0<0 To1<1 To2<1 Lo0<0 Bo0<0 Bo1<0 ]
  tran g8(.Z(w36), .I(A[3:0]));   //: @(686,-110) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g16(.Z(w14), .I(A[15:12]));   //: @(-107,-110) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  CLA g3 (.B(w37), .A(w36), .Cin(Cin), .p0(w17), .g0(w16), .S(w39));   //: @(663, 59) /sz:(162, 96) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Bo0<1 Bo1<1 Bo2<0 ]
  tran g17(.Z(w1), .I(B[11:8]));   //: @(192,-35) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  CLA g2 (.B(w27), .A(w10), .Cin(w12), .p0(w19), .g0(w18), .S(w31));   //: @(399, 60) /sz:(162, 96) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>0 Bo0<1 Bo1<1 Bo2<1 ]
  CLA g1 (.B(w1), .A(w0), .Cin(w6), .p0(w9), .g0(w20), .S(w7));   //: @(131, 56) /sz:(162, 96) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<0 Bo1<1 Bo2<0 ]
  tran g18(.Z(w27), .I(B[7:4]));   //: @(464,-35) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g10(.Z(w0), .I(A[11:8]));   //: @(157,-110) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  //: input g6 (B) @(-205,-33) /sn:0 /w:[ 0 ]
  tran g7(.Z(w37), .I(B[3:0]));   //: @(724,-35) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g9(.Z(w10), .I(A[7:4]));   //: @(415,-110) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  concat g12 (.I0(w39), .I1(w31), .I2(w7), .I3(w26), .Z(S));   //: @(884,194) /sn:0 /w:[ 1 0 1 0 0 ] /dr:0
  //: input g14 (Cin) @(991,87) /sn:0 /R:2 /w:[ 3 ]
  //: input g5 (A) @(-203,-108) /sn:0 /w:[ 9 ]
  tran g11(.Z(w2), .I(B[15:12]));   //: @(-69,-35) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: output g19 (GG) @(693,418) /sn:0 /R:3 /w:[ 1 ]
  //: output g21 (Cout) @(-258,316) /sn:0 /w:[ 1 ]
  //: output g20 (PG) @(541,416) /sn:0 /R:3 /w:[ 1 ]
  CLA g0 (.B(w2), .A(w14), .Cin(w25), .p0(w23), .g0(w22), .S(w26));   //: @(-131, 48) /sz:(162, 96) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>1 Bo0<1 Bo1<1 Bo2<1 ]
  //: joint g15 (Cin) @(971, 96) /w:[ 2 1 -1 4 ]
  //: output g13 (S) @(922,194) /sn:0 /w:[ 1 ]

endmodule

module PFA(Pi, S, Ci, B, Gi, A);
//: interface  /sz:(77, 43) /bd:[ Ti0>A(15/77) Ti1>B(44/77) Ti2>Ci(71/77) Ti3>A(14/77) Ti4>B(43/77) Ti5>Ci(70/77) Ti6>APFA(13/77) Ti7>BPFA(62/77) Ri0>CinPFA(20/43) Bo0<S(23/77) Bo1<Pi(50/77) Bo2<Gi(71/77) Bo3<S(22/77) Bo4<Pi(49/77) Bo5<Gi(70/77) Bo6<PPFA(8/77) Bo7<GFPA(20/77) Bo8<SPFA(65/77) ]
input B;    //: /sn:0 {0}(206,145)(223,145){1}
//: {2}(227,145)(269,145)(269,133)(279,133){3}
//: {4}(225,147)(225,188){5}
//: {6}(227,190)(354,190){7}
//: {8}(225,192)(225,229)(356,229){9}
output Gi;    //: /sn:0 {0}(435,225)(387,225)(387,227)(377,227){1}
input A;    //: /sn:0 {0}(205,117)(246,117){1}
//: {2}(250,117)(269,117)(269,128)(279,128){3}
//: {4}(248,119)(248,183){5}
//: {6}(250,185)(354,185){7}
//: {8}(248,187)(248,224)(356,224){9}
output Pi;    //: /sn:0 /dp:1 {0}(375,188)(422,188)(422,187)(432,187){1}
input Ci;    //: /sn:0 /dp:1 {0}(352,146)(315,146)(315,174)(204,174){1}
output S;    //: /sn:0 /dp:1 {0}(373,144)(424,144)(424,145)(433,145){1}
wire w2;    //: /sn:0 {0}(300,131)(342,131)(342,141)(352,141){1}
//: enddecls

  //: output g4 (Pi) @(429,187) /sn:0 /w:[ 1 ]
  or g8 (.I0(A), .I1(B), .Z(Pi));   //: @(365,188) /sn:0 /delay:" 3" /w:[ 7 7 0 ]
  //: output g3 (S) @(430,145) /sn:0 /w:[ 1 ]
  //: input g2 (Ci) @(202,174) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(204,145) /sn:0 /w:[ 0 ]
  //: joint g10 (A) @(248, 117) /w:[ 2 -1 1 4 ]
  xor g6 (.I0(A), .I1(B), .Z(w2));   //: @(290,131) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  xor g7 (.I0(w2), .I1(Ci), .Z(S));   //: @(363,144) /sn:0 /delay:" 4" /w:[ 1 0 0 ]
  and g9 (.I0(A), .I1(B), .Z(Gi));   //: @(367,227) /sn:0 /delay:" 3" /w:[ 9 9 1 ]
  //: joint g12 (B) @(225, 145) /w:[ 2 -1 1 4 ]
  //: output g5 (Gi) @(432,225) /sn:0 /w:[ 0 ]
  //: joint g11 (A) @(248, 185) /w:[ 6 5 -1 8 ]
  //: input g0 (A) @(203,117) /sn:0 /w:[ 0 ]
  //: joint g13 (B) @(225, 190) /w:[ 6 5 -1 8 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 /dp:1 {0}(489,352)(509,352)(509,319){1}
wire [15:0] w7;    //: /sn:0 /dp:1 {0}(397,133)(397,174){1}
wire w4;    //: /sn:0 {0}(326,233)(295,233)(295,218){1}
wire [15:0] w0;    //: /sn:0 /dp:1 {0}(536,134)(536,174){1}
wire w3;    //: /sn:0 {0}(326,286)(292,286)(292,301){1}
wire w1;    //: /sn:0 {0}(687,272)(687,250)(650,250){1}
wire [15:0] w2;    //: /sn:0 /dp:1 {0}(578,379)(578,329)(562,329)(562,319){1}
//: enddecls

  led g4 (.I(w4));   //: @(295,211) /sn:0 /w:[ 1 ] /type:0
  led g3 (.I(w6));   //: @(482,352) /sn:0 /R:1 /w:[ 0 ] /type:0
  //: dip B (w0) @(536,124) /w:[ 0 ] /st:0
  led g2 (.I(w2));   //: @(578,386) /sn:0 /R:2 /w:[ 0 ] /type:2
  //: switch g1 (w1) @(687,286) /sn:0 /R:1 /w:[ 0 ] /st:0
  //: dip A (w7) @(397,123) /w:[ 0 ] /st:18
  led g5 (.I(w3));   //: @(292,308) /sn:0 /R:2 /w:[ 1 ] /type:0
  CLA16Bits g0 (.B(w0), .A(w7), .Cin(w1), .GG(w4), .PG(w3), .S(w2), .Cout(w6));   //: @(327, 175) /sz:(322, 143) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Lo1<0 Bo0<1 Bo1<1 ]

endmodule

module CLA(A, S, B, Cin, g0, p0);
//: interface  /sz:(162, 96) /bd:[ Ti0>B[3:0](61/162) Ti1>A[3:0](24/162) Ti2>B[3:0](61/162) Ti3>A[3:0](24/162) Ri0>Cin(34/96) Ri1>Cin(34/96) Bo0<p0(130/162) Bo1<g0(87/162) Bo2<S[3:0](24/162) Bo3<p0(130/162) Bo4<g0(87/162) Bo5<S[3:0](24/162) ]
input [3:0] B;    //: /sn:0 {0}(117,75)(205,75){1}
//: {2}(206,75)(306,75){3}
//: {4}(307,75)(406,75){5}
//: {6}(407,75)(498,75){7}
//: {8}(499,75)(559,75){9}
input [3:0] A;    //: /sn:0 {0}(126,58)(175,58){1}
//: {2}(176,58)(277,58){3}
//: {4}(278,58)(378,58){5}
//: {6}(379,58)(469,58){7}
//: {8}(470,58)(557,58){9}
input Cin;    //: /sn:0 {0}(574,109)(557,109){1}
//: {2}(553,109)(526,109)(526,120){3}
//: {4}(555,111)(555,238)(538,238){5}
output p0;    //: /sn:0 {0}(483,306)(493,306)(493,292)(474,292)(474,267)(483,267)(483,257){1}
output g0;    //: /sn:0 {0}(432,303)(422,303)(422,288)(458,288)(458,257){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(639,197)(721,197){1}
wire w6;    //: /sn:0 {0}(278,123)(278,62){1}
wire w13;    //: /sn:0 {0}(407,122)(407,79){1}
wire w16;    //: /sn:0 {0}(412,164)(412,205)(413,205)(413,215){1}
wire w7;    //: /sn:0 {0}(307,123)(307,79){1}
wire w4;    //: /sn:0 {0}(201,164)(201,215){1}
wire w0;    //: /sn:0 {0}(176,122)(176,62){1}
wire w3;    //: /sn:0 {0}(174,164)(174,182)(633,182){1}
wire w22;    //: /sn:0 {0}(505,165)(505,205)(504,205)(504,215){1}
wire w20;    //: /sn:0 /dp:1 {0}(448,215)(448,112)(433,112)(433,122){1}
wire w12;    //: /sn:0 {0}(379,122)(379,62){1}
wire w18;    //: /sn:0 {0}(470,120)(470,62){1}
wire w19;    //: /sn:0 {0}(499,120)(499,79){1}
wire w10;    //: /sn:0 {0}(313,165)(313,215){1}
wire w23;    //: /sn:0 {0}(526,165)(526,205)(527,205)(527,215){1}
wire w21;    //: /sn:0 {0}(478,165)(478,212)(633,212){1}
wire w1;    //: /sn:0 {0}(206,122)(206,79){1}
wire w8;    //: /sn:0 /dp:1 {0}(250,215)(250,112)(234,112)(234,122){1}
wire w17;    //: /sn:0 {0}(433,164)(433,205)(434,205)(434,215){1}
wire w14;    //: /sn:0 /dp:1 {0}(353,215)(353,113)(334,113)(334,123){1}
wire w11;    //: /sn:0 {0}(334,165)(334,205)(335,205)(335,215){1}
wire w2;    //: /sn:0 {0}(143,237)(153,237){1}
wire w15;    //: /sn:0 {0}(386,164)(386,202)(633,202){1}
wire w5;    //: /sn:0 {0}(225,164)(225,205)(226,205)(226,215){1}
wire w9;    //: /sn:0 {0}(286,165)(286,192)(633,192){1}
//: enddecls

  //: input g4 (A) @(559,58) /sn:0 /R:2 /w:[ 9 ]
  tran g8(.Z(w0), .I(A[3]));   //: @(176,56) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  PFA g3 (.Ci(Cin), .B(w19), .A(w18), .Gi(w23), .Pi(w22), .S(w21));   //: @(455, 121) /sz:(77, 43) /sn:0 /p:[ Ti0>3 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  CLL g16 (.P3(w4), .G3(w5), .P2(w10), .G2(w11), .P1(w16), .G1(w17), .P0(w22), .G0(w23), .Cin(Cin), .C3(w8), .C2(w14), .C1(w20), .C4(w2), .PG(p0), .GG(g0));   //: @(154, 216) /sz:(383, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>5 To0<0 To1<0 To2<0 Lo0<1 Bo0<1 Bo1<1 ]
  concat g17 (.I0(w21), .I1(w15), .I2(w9), .I3(w3), .Z(S));   //: @(638,197) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  PFA g2 (.Ci(w20), .B(w13), .A(w12), .Gi(w17), .Pi(w16), .S(w15));   //: @(364, 123) /sz:(75, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  PFA g1 (.Ci(w14), .B(w7), .A(w6), .Gi(w11), .Pi(w10), .S(w9));   //: @(263, 124) /sz:(77, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  //: output g18 (S) @(718,197) /sn:0 /w:[ 1 ]
  tran g10(.Z(w19), .I(B[0]));   //: @(499,73) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g6(.Z(w12), .I(A[1]));   //: @(379,56) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g7(.Z(w6), .I(A[2]));   //: @(278,56) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: input g9 (B) @(561,75) /sn:0 /R:2 /w:[ 9 ]
  tran g12(.Z(w7), .I(B[2]));   //: @(307,73) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g5(.Z(w18), .I(A[0]));   //: @(470,56) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g11(.Z(w13), .I(B[1]));   //: @(407,73) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g14 (Cin) @(576,109) /sn:0 /R:2 /w:[ 0 ]
  //: output g19 (g0) @(429,303) /sn:0 /w:[ 0 ]
  //: output g20 (p0) @(486,306) /sn:0 /R:2 /w:[ 0 ]
  PFA g0 (.Ci(w8), .B(w1), .A(w0), .Gi(w5), .Pi(w4), .S(w3));   //: @(160, 123) /sz:(80, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  //: joint g15 (Cin) @(555, 109) /w:[ 1 -1 2 4 ]
  tran g13(.Z(w1), .I(B[3]));   //: @(206,73) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1

endmodule
