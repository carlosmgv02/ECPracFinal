//: version "1.8.7"
//: script "/home/milax/Documents/GitHub/ECPrac2/Prac2aConvo/FASE4/script.gss"


module MEM(write_data, MemRead, memWrite, read_data, Address, clk);
//: interface  /sz:(128, 174) /bd:[ Ti0>memWrite(62/128) Li0>Address[31:0](43/174) Li1>write_data[31:0](112/174) Bi0>clk(20/128) Bi1>MemRead(59/128) Ro0<read_data[31:0](27/174) ]
input [31:0] write_data;    //: /sn:0 {0}(316,166)(458,166)(458,192)(488,192){1}
output [31:0] read_data;    //: /sn:0 /dp:1 {0}(504,192)(514,192)(514,247){1}
//: {2}(516,249)(545,249){3}
//: {4}(512,249)(476,249)(476,248)(442,248){5}
input memWrite;    //: /sn:0 {0}(317,198)(353,198)(353,180)(363,180){1}
input clk;    //: /sn:0 {0}(266,135)(327,135)(327,175)(363,175){1}
supply0 w2;    //: /sn:0 {0}(338,318)(338,295)(418,295)(418,275){1}
input MemRead;    //: /sn:0 {0}(304,386)(432,386)(432,275){1}
input [31:0] Address;    //: /sn:0 {0}(379,251)(392,251)(392,250)(407,250){1}
wire w7;    //: /sn:0 {0}(384,178)(398,178){1}
//: {2}(402,178)(425,178)(425,225){3}
//: {4}(400,176)(400,153)(496,153)(496,187){5}
//: enddecls

  //: input g8 (write_data) @(314,166) /sn:0 /w:[ 0 ]
  //: input g4 (MemRead) @(302,386) /sn:0 /w:[ 0 ]
  //: input g3 (memWrite) @(315,198) /sn:0 /w:[ 0 ]
  //: output g2 (read_data) @(542,249) /sn:0 /w:[ 3 ]
  //: input g1 (Address) @(377,251) /sn:0 /w:[ 0 ]
  //: joint g6 (read_data) @(514, 249) /w:[ 2 1 4 -1 ]
  and g9 (.I0(clk), .I1(memWrite), .Z(w7));   //: @(374,178) /sn:0 /w:[ 1 1 0 ]
  //: supply0 g7 (w2) @(338,324) /sn:0 /w:[ 0 ]
  //: input g14 (clk) @(264,135) /sn:0 /w:[ 0 ]
  bufif1 g5 (.Z(read_data), .I(write_data), .E(w7));   //: @(494,192) /sn:0 /w:[ 0 1 5 ]
  //: joint g11 (w7) @(400, 178) /w:[ 2 4 1 -1 ]
  ram g0 (.A(Address), .D(read_data), .WE(!w7), .OE(!MemRead), .CS(w2));   //: @(425,249) /sn:0 /w:[ 1 5 3 1 1 ]

endmodule

module ALUCtrl(ALUOp, ALUCtrl, funct);
//: interface  /sz:(134, 106) /bd:[ Li0>funct[5:0](51/106) Li1>ALUOp[1:0](17/106) Ro0<ALUCtrl[3:0](24/106) ]
output [3:0] ALUCtrl;    //: /sn:0 /dp:1 {0}(1002,416)(1057,416)(1057,423)(1106,423){1}
supply0 [3:0] w4;    //: /sn:0 {0}(839,369)(839,398)(973,398){1}
supply0 w3;    //: /sn:0 {0}(610,456)(610,444){1}
input [1:0] ALUOp;    //: /sn:0 {0}(314,545)(989,545)(989,439){1}
input [5:0] funct;    //: /sn:0 {0}(407,426)(526,426)(526,419)(592,419){1}
wire [3:0] w0;    //: /sn:0 {0}(723,451)(881,451)(881,422)(973,422){1}
wire [3:0] w1;    //: /sn:0 {0}(627,417)(805,417)(805,410)(973,410){1}
wire [3:0] w2;    //: /sn:0 {0}(822,482)(963,482)(963,434)(973,434){1}
//: enddecls

  //: input g4 (ALUOp) @(312,545) /sn:0 /w:[ 0 ]
  //: output g8 (ALUCtrl) @(1103,423) /sn:0 /w:[ 1 ]
  mux g3 (.I0(w2), .I1(w0), .I2(w1), .I3(w4), .S(ALUOp), .Z(ALUCtrl));   //: @(989,416) /sn:0 /R:1 /w:[ 1 1 1 1 1 0 ] /ss:0 /do:0
  //: input g2 (funct) @(405,426) /sn:0 /w:[ 0 ]
  //: supply0 g1 (w3) @(610,462) /sn:0 /w:[ 0 ]
  //: dip g6 (w0) @(685,451) /sn:0 /R:1 /w:[ 0 ] /st:6
  //: supply0 g7 (w4) @(839,363) /sn:0 /R:2 /w:[ 0 ]
  //: dip g5 (w2) @(784,482) /sn:0 /R:1 /w:[ 0 ] /st:2
  rom g0 (.A(funct), .D(w1), .OE(w3));   //: @(610,418) /sn:0 /w:[ 1 0 1 ]

endmodule

module CSA(B, A, Cin, S, Cout);
//: interface  /sz:(127, 64) /bd:[ Ti0>A[3:0](9/127) Ti1>B[3:0](30/127) Ti2>Cin(74/127) To0<Cout(96/127) To1<S[3:0](48/127) ]
input [3:0] B;    //: /sn:0 /dp:5 {0}(572,36)(490,36){1}
//: {2}(489,36)(458,36)(458,36)(372,36){3}
//: {4}(371,36)(265,36)(265,44)(256,44){5}
//: {6}(255,44)(144,44){7}
//: {8}(143,44)(42,44){9}
input [3:0] A;    //: /sn:0 {0}(43,23)(173,23){1}
//: {2}(174,23)(278,23)(278,7)(285,7){3}
//: {4}(286,7)(294,7)(294,23)(404,23){5}
//: {6}(405,23)(521,23){7}
//: {8}(522,23)(565,23){9}
supply0 w10;    //: /sn:0 {0}(527,105)(591,105)(591,106)(601,106){1}
input Cin;    //: /sn:0 {0}(613,304)(464,304)(464,313){1}
//: {2}(462,315)(346,315)(346,318){3}
//: {4}(344,320)(235,320)(235,321)(225,321){5}
//: {6}(221,321)(104,321)(104,340){7}
//: {8}(106,342)(118,342)(118,343)(130,343){9}
//: {10}(102,342)(39,342)(39,133)(57,133)(57,143){11}
//: {12}(223,323)(223,338)(246,338){13}
//: {14}(346,322)(346,335)(368,335){15}
//: {16}(464,317)(464,335)(490,335){17}
output Cout;    //: /sn:0 {0}(1,165)(32,165)(32,166)(44,166){1}
supply1 w11;    //: /sn:0 {0}(644,230)(597,230)(597,231)(552,231){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(570,405)(604,405){1}
wire w13;    //: /sn:0 /dp:1 {0}(259,134)(259,322){1}
wire w50;    //: /sn:0 {0}(391,348)(391,410)(564,410){1}
wire w4;    //: /sn:0 {0}(133,139)(133,156)(73,156){1}
wire w25;    //: /sn:0 {0}(301,236)(317,236)(317,286)(349,286)(349,298)(379,298)(379,268){1}
wire w0;    //: /sn:0 {0}(275,199)(275,184)(313,184)(313,55)(288,55){1}
//: {2}(286,53)(286,11){3}
//: {4}(286,57)(286,79){5}
wire w22;    //: /sn:0 {0}(139,201)(139,187)(154,187)(154,60)(146,60){1}
//: {2}(144,58)(144,48){3}
//: {4}(144,62)(144,76){5}
wire w36;    //: /sn:0 {0}(528,193)(528,184)(542,184)(542,58)(525,58){1}
//: {2}(523,56)(523,31)(522,31)(522,27){3}
//: {4}(523,60)(523,67)(501,67)(501,72){5}
wire w20;    //: /sn:0 {0}(187,235)(193,235)(193,292)(237,292)(237,278){1}
wire w30;    //: /sn:0 {0}(428,230)(443,230)(443,291)(495,291)(495,273){1}
wire w37;    //: /sn:0 /dp:1 {0}(490,40)(490,46)(489,46)(489,56){1}
//: {2}(491,58)(512,58)(512,181)(500,181)(500,193){3}
//: {4}(489,60)(489,67)(467,67)(467,72){5}
wire w19;    //: /sn:0 {0}(510,142)(510,163)(429,163)(429,103)(419,103){1}
wire w23;    //: /sn:0 {0}(162,274)(162,317)(163,317)(163,327){1}
wire w54;    //: /sn:0 {0}(513,348)(513,420)(564,420){1}
wire w21;    //: /sn:0 {0}(165,201)(165,186)(185,186)(185,63)(175,63){1}
//: {2}(173,61)(173,36)(174,36)(174,27){3}
//: {4}(173,65)(173,76){5}
wire w24;    //: /sn:0 {0}(153,356)(153,390)(564,390){1}
wire w31;    //: /sn:0 {0}(403,197)(403,181)(422,181)(422,56)(407,56){1}
//: {2}(405,54)(405,27){3}
//: {4}(405,58)(405,66)(396,66)(396,73){5}
wire w1;    //: /sn:0 {0}(357,141)(357,302)(381,302)(381,319){1}
wire w32;    //: /sn:0 /dp:1 {0}(372,40)(372,56){1}
//: {2}(374,58)(387,58)(387,184)(371,184)(371,197){3}
//: {4}(372,60)(372,67)(363,67)(363,73){5}
wire w46;    //: /sn:0 {0}(269,351)(269,400)(564,400){1}
wire w8;    //: /sn:0 {0}(301,105)(322,105)(322,165)(403,165)(403,141){1}
wire w27;    //: /sn:0 {0}(245,199)(245,188)(269,188)(269,65)(252,65){1}
//: {2}(250,63)(250,56)(256,56)(256,48){3}
//: {4}(250,67)(250,79){5}
wire w28;    //: /sn:0 {0}(272,278)(272,301)(279,301)(279,322){1}
wire w33;    //: /sn:0 {0}(408,268)(408,309)(401,309)(401,319){1}
wire w41;    //: /sn:0 /dp:1 {0}(73,176)(87,176)(87,301)(134,301)(134,274){1}
wire w2;    //: /sn:0 {0}(287,134)(287,155)(222,155)(222,105)(194,105){1}
wire w38;    //: /sn:0 {0}(525,273)(525,309)(523,309)(523,319){1}
wire w9;    //: /sn:0 /dp:1 {0}(143,327)(143,312)(158,312)(158,139){1}
wire w51;    //: /sn:0 /dp:1 {0}(503,319)(503,311)(476,311)(476,142){1}
//: enddecls

  concat g44 (.I0(w54), .I1(w50), .I2(w46), .I3(w24), .Z(S));   //: @(569,405) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  FA g4 (.B(w22), .A(w21), .Cin(w20), .Cout(w41), .S(w23));   //: @(120, 202) /sz:(66, 71) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Bo0<1 Bo1<0 ]
  mux g8 (.I0(w4), .I1(w41), .S(Cin), .Z(Cout));   //: @(57,166) /sn:0 /R:3 /delay:" 2 2" /w:[ 1 0 11 1 ] /ss:0 /do:0
  tran g16(.Z(w0), .I(A[2]));   //: @(286,5) /sn:0 /R:1 /w:[ 3 3 4 ] /ss:1
  FA g3 (.B(w37), .A(w36), .Cin(w10), .Cout(w19), .S(w51));   //: @(447, 73) /sz:(79, 68) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Bo0<0 Bo1<1 ]
  tran g26(.Z(w21), .I(A[3]));   //: @(174,21) /sn:0 /R:1 /w:[ 3 1 2 ] /ss:1
  //: joint g17 (w32) @(372, 58) /w:[ 2 1 -1 4 ]
  FA g2 (.B(w32), .A(w31), .Cin(w19), .Cout(w8), .S(w1));   //: @(340, 74) /sz:(79, 66) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>1 Bo0<1 Bo1<0 ]
  //: joint g23 (Cin) @(346, 320) /w:[ -1 3 4 14 ]
  //: input g30 (B) @(40,44) /sn:0 /w:[ 9 ]
  //: joint g24 (Cin) @(464, 315) /w:[ -1 1 2 16 ]
  FA g1 (.B(w27), .A(w0), .Cin(w8), .Cout(w2), .S(w13));   //: @(235, 80) /sz:(65, 53) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Bo0<0 Bo1<0 ]
  tran g29(.Z(w36), .I(A[0]));   //: @(522,21) /sn:0 /R:1 /w:[ 3 7 8 ] /ss:1
  //: joint g18 (w31) @(405, 56) /w:[ 1 2 -1 4 ]
  mux g10 (.I0(w13), .I1(w28), .S(Cin), .Z(w46));   //: @(269,338) /sn:0 /delay:" 2 2" /w:[ 1 1 13 0 ] /ss:0 /do:0
  //: input g25 (A) @(41,23) /sn:0 /w:[ 0 ]
  FA g6 (.B(w32), .A(w31), .Cin(w30), .Cout(w25), .S(w33));   //: @(351, 198) /sz:(76, 69) /sn:0 /p:[ Ti0>3 Ti1>0 Ri0>0 Bo0<1 Bo1<0 ]
  //: input g35 (Cin) @(615,304) /sn:0 /R:2 /w:[ 0 ]
  FA g7 (.B(w37), .A(w36), .Cin(w11), .Cout(w30), .S(w38));   //: @(481, 194) /sz:(71, 78) /sn:0 /p:[ Ti0>3 Ti1>0 Ri0>1 Bo0<1 Bo1<0 ]
  mux g9 (.I0(w9), .I1(w23), .S(Cin), .Z(w24));   //: @(153,343) /sn:0 /delay:" 2 2" /w:[ 0 1 9 0 ] /ss:0 /do:0
  //: joint g31 (w27) @(250, 65) /w:[ 1 2 -1 4 ]
  //: joint g22 (Cin) @(223, 321) /w:[ 5 -1 6 12 ]
  //: supply0 g36 (w10) @(607,106) /sn:0 /R:1 /w:[ 1 ]
  tran g33(.Z(w32), .I(B[1]));   //: @(372,34) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  mux g12 (.I0(w51), .I1(w38), .S(Cin), .Z(w54));   //: @(513,335) /sn:0 /delay:" 2 2" /w:[ 0 1 17 0 ] /ss:0 /do:0
  tran g28(.Z(w31), .I(A[1]));   //: @(405,21) /sn:0 /R:1 /w:[ 3 5 6 ] /ss:1
  tran g34(.Z(w37), .I(B[0]));   //: @(490,34) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  FA g5 (.B(w27), .A(w0), .Cin(w25), .Cout(w20), .S(w28));   //: @(224, 200) /sz:(77, 77) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Bo0<1 Bo1<0 ]
  mux g11 (.I0(w1), .I1(w33), .S(Cin), .Z(w50));   //: @(391,335) /sn:0 /delay:" 2 2" /w:[ 1 1 15 0 ] /ss:0 /do:0
  //: joint g14 (w21) @(173, 63) /w:[ 1 2 -1 4 ]
  //: joint g21 (Cin) @(104, 342) /w:[ 8 7 10 -1 ]
  //: joint g19 (w37) @(489, 58) /w:[ 2 1 -1 4 ]
  //: joint g20 (w36) @(523, 58) /w:[ 1 2 -1 4 ]
  tran g32(.Z(w22), .I(B[3]));   //: @(144,42) /sn:0 /R:1 /w:[ 3 8 7 ] /ss:1
  //: output g38 (S) @(601,405) /sn:0 /w:[ 1 ]
  tran g15(.Z(w27), .I(B[2]));   //: @(256,42) /sn:0 /R:1 /w:[ 3 6 5 ] /ss:1
  //: supply1 g43 (w11) @(644,241) /sn:0 /R:3 /w:[ 0 ]
  FA g0 (.B(w22), .A(w21), .Cin(w2), .Cout(w4), .S(w9));   //: @(119, 77) /sz:(75, 61) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>1 Bo0<0 Bo1<1 ]
  //: joint g27 (w0) @(286, 55) /w:[ 1 2 -1 4 ]
  //: output g37 (Cout) @(4,165) /sn:0 /R:2 /w:[ 0 ]
  //: joint g13 (w22) @(144, 60) /w:[ 1 2 -1 4 ]

endmodule

module CLA32(Cout, B, A, S, Cin);
//: interface  /sz:(136, 114) /bd:[ Ti0>A[31:0](32/136) Ti1>B[31:0](92/136) Ri0>Cin(60/114) Lo0<Cout(62/114) Bo0<S[31:0](68/136) ]
input [31:0] B;    //: /sn:0 {0}(1071,151)(887,151){1}
//: {2}(886,151)(497,151){3}
//: {4}(496,151)(247,151){5}
input [31:0] A;    //: /sn:0 {0}(1065,95)(750,95){1}
//: {2}(749,95)(350,95){3}
//: {4}(349,95)(229,95){5}
input Cin;    //: /sn:0 {0}(950,392)(1001,392)(1001,381)(1011,381)(1011,395)(1069,395){1}
output Cout;    //: /sn:0 {0}(480,507)(464,507)(464,446){1}
output [31:0] S;    //: /sn:0 /dp:1 {0}(884,601)(916,601)(916,593)(926,593){1}
wire [15:0] w13;    //: /sn:0 /dp:1 {0}(878,606)(799,606)(799,507)(857,507)(857,451){1}
wire [15:0] w6;    //: /sn:0 {0}(753,321)(753,107)(750,107)(750,99){1}
wire w4;    //: /sn:0 /dp:1 {0}(262,467)(262,413)(281,413){1}
wire [15:0] w0;    //: /sn:0 {0}(352,301)(352,107)(350,107)(350,99){1}
wire [15:0] w3;    //: /sn:0 {0}(870,321)(870,305)(887,305)(887,155){1}
wire w12;    //: /sn:0 {0}(605,377)(659,377)(659,482)(744,482)(744,451){1}
wire [15:0] w1;    //: /sn:0 {0}(491,301)(491,163)(497,163)(497,155){1}
wire w2;    //: /sn:0 /dp:1 {0}(257,339)(257,360)(281,360){1}
wire [15:0] w5;    //: /sn:0 /dp:1 {0}(878,596)(517,596)(517,446){1}
//: enddecls

  //: output g8 (Cout) @(477,507) /sn:0 /w:[ 0 ]
  tran g4(.Z(w3), .I(B[15:0]));   //: @(887,149) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  //: input g3 (B) @(1073,151) /sn:0 /R:2 /w:[ 0 ]
  //: input g2 (A) @(1067,95) /sn:0 /R:2 /w:[ 0 ]
  CSA16bits g1 (.A(w6), .B(w3), .Cin(Cin), .S(w13), .Cout(w12));   //: @(692, 322) /sz:(257, 128) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Bo0<1 Bo1<1 ]
  //: output g10 (S) @(923,593) /sn:0 /w:[ 1 ]
  tran g6(.Z(w1), .I(B[31:16]));   //: @(497,149) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  concat g9 (.I0(w13), .I1(w5), .Z(S));   //: @(883,601) /sn:0 /w:[ 0 0 0 ] /dr:0
  tran g7(.Z(w0), .I(A[31:16]));   //: @(350,93) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  led g12 (.I(w4));   //: @(262,474) /sn:0 /R:2 /w:[ 0 ] /type:0
  led g11 (.I(w2));   //: @(257,332) /sn:0 /w:[ 0 ] /type:0
  tran g5(.Z(w6), .I(A[15:0]));   //: @(750,93) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  //: input g15 (Cin) @(1071,395) /sn:0 /R:2 /w:[ 1 ]
  CLA16Bits g0 (.B(w1), .A(w0), .Cin(w12), .GG(w2), .PG(w4), .S(w5), .Cout(Cout));   //: @(282, 302) /sz:(322, 143) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Lo1<1 Bo0<1 Bo1<1 ]

endmodule

module ctrl(RegDst, ALUSrc, op, MemRead, Jump, cmpseti, MemtoReg, Branch, RegWrite, funct, MemWrite, ALUCtrl);
//: interface  /sz:(171, 204) /bd:[ Li0>op[5:0](34/204) Li1>funct[5:0](149/204) Ro0<RegDst(16/204) Ro1<Jump(31/204) Ro2<Branch(49/204) Ro3<MemRead(67/204) Ro4<ALUCtrl[3:0](111/204) Ro5<MemtoReg(88/204) Ro6<MemWrite(129/204) Ro7<ALUSrc(155/204) Ro8<RegWrite(177/204) ]
output cmpseti;    //: /sn:0 /dp:1 {0}(849,160)(942,160){1}
output Branch;    //: /sn:0 {0}(849,215)(978,215){1}
output [3:0] ALUCtrl;    //: /sn:0 /dp:1 {0}(849,387)(857,387)(857,388)(994,388){1}
supply0 w3;    //: /sn:0 {0}(726,251)(726,193)(748,193)(748,183){1}
output MemWrite;    //: /sn:0 {0}(849,436)(857,436)(857,437)(982,437){1}
output [1:0] ALUSrc;    //: /sn:0 {0}(849,470)(916,470)(916,471)(1005,471){1}
output RegDst;    //: /sn:0 {0}(849,181)(975,181){1}
output RegWrite;    //: /sn:0 {0}(849,502)(857,502)(857,501)(1002,501){1}
output MemtoReg;    //: /sn:0 {0}(850,329)(858,329)(858,337)(980,337){1}
output MemRead;    //: /sn:0 {0}(849,286)(857,286)(857,291)(983,291){1}
input [5:0] funct;    //: /sn:0 {0}(559,199)(423,199){1}
input [5:0] op;    //: /sn:0 {0}(429,179)(444,179){1}
//: {2}(445,179)(471,179){3}
//: {4}(472,179)(488,179){5}
//: {6}(489,179)(505,179){7}
//: {8}(506,179)(524,179){9}
//: {10}(525,179)(540,179){11}
//: {12}(541,179)(559,179){13}
output Jump;    //: /sn:0 {0}(849,252)(857,252)(857,255)(980,255){1}
wire [1:0] w6;    //: /sn:0 /dp:1 {0}(642,309)(642,280)(650,280)(650,204)(671,204){1}
wire w7;    //: /sn:0 {0}(563,264)(575,264)(575,212){1}
wire w4;    //: /sn:0 {0}(525,183)(525,257)(542,257){1}
wire [7:0] w0;    //: /sn:0 {0}(730,158)(687,158)(687,209)(677,209){1}
wire w10;    //: /sn:0 {0}(542,272)(472,272)(472,183){1}
wire [15:0] w1;    //: /sn:0 /dp:1 {0}(765,156)(810,156){1}
//: {2}(814,156)(845,156)(845,159){3}
//: {4}(845,160)(845,180){5}
//: {6}(845,181)(845,214){7}
//: {8}(845,215)(845,251){9}
//: {10}(845,252)(845,285){11}
//: {12}(845,286)(845,306)(846,306)(846,328){13}
//: {14}(846,329)(846,376)(845,376)(845,386){15}
//: {16}(845,387)(845,435){17}
//: {18}(845,436)(845,469){19}
//: {20}(845,470)(845,501){21}
//: {22}(845,502)(845,655){23}
//: {24}(812,154)(812,144)(814,144)(814,70){25}
wire w8;    //: /sn:0 {0}(542,262)(506,262)(506,183){1}
wire w2;    //: /sn:0 {0}(541,183)(541,252)(542,252){1}
wire w11;    //: /sn:0 {0}(542,277)(445,277)(445,183){1}
wire [5:0] w5;    //: /sn:0 {0}(671,214)(612,214)(612,189)(588,189){1}
wire w9;    //: /sn:0 {0}(542,267)(489,267)(489,183){1}
//: enddecls

  tran g8(.Z(Jump), .I(w1[12]));   //: @(843,252) /sn:0 /R:2 /w:[ 0 10 9 ] /ss:1
  tran g4(.Z(RegDst), .I(w1[14]));   //: @(843,181) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  //: output g3 (RegDst) @(972,181) /sn:0 /w:[ 1 ]
  tran g16(.Z(MemWrite), .I(w1[3]));   //: @(843,436) /sn:0 /R:2 /w:[ 0 18 17 ] /ss:1
  //: output g17 (ALUSrc) @(1002,471) /sn:0 /w:[ 1 ]
  tran g26(.Z(w8), .I(op[3]));   //: @(506,177) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: input g2 (op) @(427,179) /sn:0 /w:[ 0 ]
  or g23 (.I0(w2), .I1(w4), .I2(w8), .I3(w9), .I4(w10), .I5(w11), .Z(w7));   //: @(553,264) /sn:0 /w:[ 1 1 0 0 0 0 0 ]
  concat g30 (.I0(w5), .I1(w6), .Z(w0));   //: @(676,209) /sn:0 /w:[ 0 1 1 ] /dr:0
  //: supply0 g1 (w3) @(726,257) /sn:0 /w:[ 0 ]
  tran g24(.Z(w2), .I(op[5]));   //: @(541,177) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  tran g29(.Z(w11), .I(op[0]));   //: @(445,177) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g18(.Z(ALUSrc), .I(w1[2:1]));   //: @(843,470) /sn:0 /R:2 /w:[ 0 20 19 ] /ss:1
  tran g10(.Z(MemRead), .I(w1[11]));   //: @(843,286) /sn:0 /R:2 /w:[ 0 12 11 ] /ss:1
  tran g25(.Z(w4), .I(op[4]));   //: @(525,177) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  tran g6(.Z(Branch), .I(w1[13]));   //: @(843,215) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  //: output g9 (MemRead) @(980,291) /sn:0 /w:[ 1 ]
  //: output g7 (Jump) @(977,255) /sn:0 /w:[ 1 ]
  tran g35(.Z(cmpseti), .I(w1[15]));   //: @(843,160) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  mux g22 (.I0(funct), .I1(op), .S(w7), .Z(w5));   //: @(575,189) /sn:0 /R:1 /w:[ 0 13 1 1 ] /ss:0 /do:0
  //: dip g31 (w6) @(642,320) /sn:0 /R:2 /w:[ 0 ] /st:0
  //: joint g33 (w1) @(812, 156) /w:[ 2 24 1 -1 ]
  tran g12(.Z(MemtoReg), .I(w1[10]));   //: @(844,329) /sn:0 /R:2 /w:[ 0 14 13 ] /ss:1
  tran g28(.Z(w10), .I(op[1]));   //: @(472,177) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: output g34 (cmpseti) @(939,160) /sn:0 /w:[ 1 ]
  //: output g11 (MemtoReg) @(977,337) /sn:0 /w:[ 1 ]
  //: output g5 (Branch) @(975,215) /sn:0 /w:[ 1 ]
  tran g14(.Z(ALUCtrl), .I(w1[9:6]));   //: @(843,387) /sn:0 /R:2 /w:[ 0 16 15 ] /ss:1
  //: output g19 (RegWrite) @(999,501) /sn:0 /w:[ 1 ]
  //: input g21 (funct) @(421,199) /sn:0 /w:[ 1 ]
  led g32 (.I(w1));   //: @(814,63) /sn:0 /w:[ 25 ] /type:1
  tran g20(.Z(RegWrite), .I(w1[0]));   //: @(843,502) /sn:0 /R:2 /w:[ 0 22 21 ] /ss:1
  rom g0 (.A(w0), .D(w1), .OE(w3));   //: @(748,157) /sn:0 /w:[ 0 0 1 ]
  //: output g15 (MemWrite) @(979,437) /sn:0 /w:[ 1 ]
  tran g27(.Z(w9), .I(op[2]));   //: @(489,177) /sn:0 /R:1 /anc:1 /w:[ 1 5 6 ] /ss:1
  //: output g13 (ALUCtrl) @(991,388) /sn:0 /w:[ 1 ]

endmodule

module READ(Read_register_2, Read_data_2, Pop, Write_register, mux_RegDst, Read_register_1, clk, Write_data, Sign_ext_out, Sign_ext_in, clr, Read_data_1, RegWrite);
//: interface  /sz:(255, 283) /bd:[ Ti0>Pop(49/255) Ti1>RegWrite(135/255) Li0>Read_register_1[4:0](51/283) Li1>Read_register_2[4:0](102/283) Li2>Write_register[4:0](151/283) Li3>mux_RegDst(180/283) Li4>Sign_ext_in[15:0](237/283) Bi0>clk(87/255) Bi1>clr(144/255) Bi2>Write_data[31:0](20/255) Ro0<Read_data_1[31:0](53/283) Ro1<Read_data_2[31:0](162/283) Ro2<Sign_ext_out[31:0](250/283) ]
input Pop;    //: /sn:0 {0}(568,-9)(440,-9)(440,34){1}
output [31:0] Read_data_1;    //: /sn:0 /dp:1 {0}(483,82)(616,82)(616,83)(626,83){1}
input [4:0] Write_register;    //: /sn:0 {0}(66,173)(150,173)(150,133)(170,133){1}
input [4:0] Read_register_1;    //: /sn:0 /dp:1 {0}(83,67)(334,67){1}
input [4:0] Read_register_2;    //: /sn:0 /dp:1 {0}(89,133)(118,133){1}
//: {2}(120,131)(120,107)(334,107){3}
//: {4}(120,135)(120,153)(170,153){5}
output [31:0] Read_data_2;    //: /sn:0 /dp:1 {0}(483,174)(561,174)(561,165)(571,165){1}
input [31:0] Write_data;    //: /sn:0 /dp:1 {0}(94,235)(242,235)(242,183)(334,183){1}
input RegWrite;    //: /sn:0 {0}(7,290)(375,290)(375,218){1}
input clr;    //: /sn:0 {0}(259,-43)(401,-43)(401,34){1}
input mux_RegDst;    //: /sn:0 {0}(94,210)(186,210)(186,166){1}
output [31:0] Sign_ext_out;    //: /sn:0 /dp:1 {0}(420,408)(597,408)(597,407)(618,407){1}
input clk;    //: /sn:0 {0}(462,356)(462,287)(455,287)(455,256)(445,256){1}
//: {2}(443,254)(443,218){3}
//: {4}(443,258)(443,266){5}
input [15:0] Sign_ext_in;    //: /sn:0 {0}(62,403)(315,403){1}
wire [4:0] w3;    //: /sn:0 /dp:1 {0}(199,143)(334,143){1}
//: enddecls

  BRegs32x32 g4 (.Pop(Pop), .clr(clr), .Read1(Read_register_1), .Read2(Read_register_2), .Write(w3), .WriteData(Write_data), .clk(clk), .RegWrite(RegWrite), .Data1(Read_data_1), .Data2(Read_data_2));   //: @(335, 35) /sz:(147, 182) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Li1>3 Li2>1 Li3>1 Bi0>3 Bi1>1 Ro0<0 Ro1<0 ]
  //: joint g8 (clk) @(443, 256) /w:[ 1 2 -1 4 ]
  //: input g3 (Read_register_2) @(87,133) /sn:0 /w:[ 0 ]
  //: output g16 (Read_data_2) @(568,165) /sn:0 /w:[ 1 ]
  //: input g17 (Pop) @(570,-9) /sn:0 /R:2 /w:[ 0 ]
  //: input g2 (Write_register) @(64,173) /sn:0 /w:[ 0 ]
  //: input g1 (mux_RegDst) @(92,210) /sn:0 /w:[ 0 ]
  signextend g10 (.In(Sign_ext_in), .Out(Sign_ext_out));   //: @(316, 373) /sz:(103, 81) /sn:0 /p:[ Li0>1 Ro0<0 ]
  //: input g6 (Read_register_1) @(81,67) /sn:0 /w:[ 0 ]
  //: input g9 (clk) @(462,358) /sn:0 /R:1 /w:[ 0 ]
  //: input g7 (Write_data) @(92,235) /sn:0 /w:[ 0 ]
  //: output g12 (Sign_ext_out) @(615,407) /sn:0 /w:[ 1 ]
  //: joint g5 (Read_register_2) @(120, 133) /w:[ -1 2 1 4 ]
  //: input g11 (Sign_ext_in) @(60,403) /sn:0 /w:[ 0 ]
  //: input g14 (clr) @(257,-43) /sn:0 /w:[ 0 ]
  mux g0 (.I0(Read_register_2), .I1(Write_register), .S(mux_RegDst), .Z(w3));   //: @(186,143) /sn:0 /R:1 /w:[ 5 1 1 0 ] /ss:0 /do:0
  //: output g15 (Read_data_1) @(623,83) /sn:0 /w:[ 1 ]
  //: input g13 (RegWrite) @(5,290) /sn:0 /w:[ 0 ]

endmodule

module CLL(G3, P1, G1, G0, Cin, G2, P2, PG, C2, C4, C1, P3, P0, GG, C3);
//: interface  /sz:(974, 86) /bd:[ Ti0>P3(120/974) Ti1>G3(182/974) Ti2>P2(402/974) Ti3>G2(457/974) Ti4>P1(657/974) Ti5>G1(710/974) Ti6>P0(887/974) Ti7>G0(946/974) Ri0>Cin(57/86) To0<C3(242/974) To1<C2(505/974) To2<C1(746/974) Lo0<C4(45/86) Bo0<PG(685/974) Bo1<GG(837/974) ]
input G2;    //: /sn:0 {0}(297,703)(267,703){1}
//: {2}(265,701)(265,518){3}
//: {4}(267,516)(362,516){5}
//: {6}(263,516)(167,516){7}
//: {8}(265,705)(265,851)(299,851){9}
output GG;    //: /sn:0 {0}(427,807)(398,807){1}
input P1;    //: /sn:0 {0}(300,782)(243,782)(243,742){1}
//: {2}(245,740)(299,740){3}
//: {4}(243,738)(243,634){5}
//: {6}(245,632)(298,632){7}
//: {8}(243,630)(243,590){9}
//: {10}(245,588)(298,588){11}
//: {12}(243,586)(243,523)(216,523)(216,506){13}
//: {14}(218,504)(286,504){15}
//: {16}(216,502)(216,474){17}
//: {18}(218,472)(287,472){19}
//: {20}(216,470)(216,410){21}
//: {22}(218,408)(286,408){23}
//: {24}(216,406)(216,374){25}
//: {26}(218,372)(287,372){27}
//: {28}(214,372)(166,372){29}
output C3;    //: /sn:0 {0}(408,508)(383,508){1}
output PG;    //: /sn:0 /dp:1 {0}(320,742)(364,742){1}
input G0;    //: /sn:0 /dp:1 {0}(334,261)(261,261)(261,294)(211,294){1}
//: {2}(207,294)(177,294)(177,309)(167,309){3}
//: {4}(209,296)(209,411){5}
//: {6}(211,413)(286,413){7}
//: {8}(209,415)(209,497){9}
//: {10}(211,499)(286,499){11}
//: {12}(209,501)(209,625){13}
//: {14}(211,627)(298,627){15}
//: {16}(209,629)(209,777)(300,777){17}
output C4;    //: /sn:0 {0}(438,655)(403,655){1}
output C2;    //: /sn:0 {0}(401,385)(369,385){1}
input Cin;    //: /sn:0 /dp:7 {0}(287,362)(232,362){1}
//: {2}(230,360)(230,287){3}
//: {4}(230,283)(230,258)(235,258){5}
//: {6}(228,285)(167,285){7}
//: {8}(230,364)(230,460){9}
//: {10}(232,462)(287,462){11}
//: {12}(230,464)(230,578)(298,578){13}
input P3;    //: /sn:0 /dp:1 {0}(299,745)(260,745){1}
//: {2}(258,743)(258,710){3}
//: {4}(260,708)(297,708){5}
//: {6}(258,706)(258,680){7}
//: {8}(260,678)(298,678){9}
//: {10}(258,676)(258,644){11}
//: {12}(260,642)(298,642){13}
//: {14}(258,640)(258,600){15}
//: {16}(260,598)(298,598){17}
//: {18}(256,598)(170,598)(170,598)(167,598){19}
//: {20}(258,747)(258,790){21}
//: {22}(260,792)(300,792){23}
//: {24}(258,794)(258,824){25}
//: {26}(260,826)(300,826){27}
//: {28}(258,828)(258,856)(299,856){29}
input G1;    //: /sn:0 {0}(166,385)(200,385){1}
//: {2}(204,385)(348,385){3}
//: {4}(202,387)(202,511){5}
//: {6}(204,513)(279,513)(279,536)(289,536){7}
//: {8}(202,515)(202,666){9}
//: {10}(204,668)(298,668){11}
//: {12}(202,670)(202,816)(300,816){13}
input G3;    //: /sn:0 /dp:1 {0}(382,655)(224,655){1}
//: {2}(220,655)(166,655){3}
//: {4}(222,657)(222,805)(377,805){5}
output C1;    //: /sn:0 /dp:1 {0}(355,259)(399,259){1}
input P0;    //: /sn:0 {0}(287,467)(238,467){1}
//: {2}(236,465)(236,369){3}
//: {4}(238,367)(287,367){5}
//: {6}(234,367)(221,367)(221,236){7}
//: {8}(223,234)(229,234)(229,253)(235,253){9}
//: {10}(219,234)(180,234)(180,234)(166,234){11}
//: {12}(236,469)(236,581){13}
//: {14}(238,583)(298,583){15}
//: {16}(236,585)(236,735)(299,735){17}
input P2;    //: /sn:0 {0}(299,750)(275,750){1}
//: {2}(273,748)(273,675){3}
//: {4}(275,673)(298,673){5}
//: {6}(271,673)(250,673)(250,639){7}
//: {8}(252,637)(298,637){9}
//: {10}(250,635)(250,595){11}
//: {12}(252,593)(298,593){13}
//: {14}(250,591)(250,511){15}
//: {16}(252,509)(286,509){17}
//: {18}(248,509)(227,509){19}
//: {20}(225,507)(225,479){21}
//: {22}(227,477)(287,477){23}
//: {24}(223,477)(168,477){25}
//: {26}(225,511)(225,541)(289,541){27}
//: {28}(273,752)(273,785){29}
//: {30}(275,787)(300,787){31}
//: {32}(273,789)(273,821)(300,821){33}
wire w6;    //: /sn:0 {0}(320,854)(367,854)(367,815)(377,815){1}
wire w4;    //: /sn:0 {0}(321,784)(367,784)(367,800)(377,800){1}
wire w39;    //: /sn:0 /dp:1 {0}(318,706)(345,706)(345,665)(382,665){1}
wire w3;    //: /sn:0 {0}(307,411)(338,411)(338,390)(348,390){1}
wire D8;    //: /sn:0 {0}(308,367)(338,367)(338,380)(348,380){1}
wire w42;    //: /sn:0 /dp:1 {0}(319,588)(346,588)(346,645)(382,645){1}
wire w18;    //: /sn:0 /dp:1 {0}(307,504)(317,504)(317,506)(362,506){1}
wire w8;    //: /sn:0 {0}(377,810)(359,810)(359,821)(321,821){1}
wire w44;    //: /sn:0 {0}(362,511)(320,511)(320,539)(310,539){1}
wire w45;    //: /sn:0 /dp:1 {0}(308,469)(321,469)(321,501)(362,501){1}
wire w2;    //: /sn:0 /dp:1 {0}(256,256)(334,256){1}
wire w15;    //: /sn:0 /dp:1 {0}(319,634)(340,634)(340,650)(382,650){1}
wire w40;    //: /sn:0 /dp:1 {0}(319,673)(339,673)(339,660)(382,660){1}
//: enddecls

  and g44 (.I0(G1), .I1(P2), .I2(P3), .Z(w40));   //: @(309,673) /sn:0 /delay:" 3" /w:[ 11 5 9 0 ]
  //: input g8 (G3) @(164,655) /sn:0 /w:[ 3 ]
  //: input g4 (P1) @(164,372) /sn:0 /w:[ 29 ]
  //: joint g47 (P3) @(258, 642) /w:[ 12 14 -1 11 ]
  //: joint g16 (Cin) @(230, 285) /w:[ -1 4 6 3 ]
  //: input g3 (G1) @(164,385) /sn:0 /w:[ 0 ]
  //: joint g17 (P0) @(221, 234) /w:[ 8 -1 10 7 ]
  and g26 (.I0(G0), .I1(P1), .I2(P2), .Z(w18));   //: @(297,504) /sn:0 /delay:" 3" /w:[ 11 15 17 0 ]
  //: input g2 (G0) @(165,309) /sn:0 /w:[ 3 ]
  //: joint g23 (Cin) @(230, 362) /w:[ 1 2 -1 8 ]
  and g30 (.I0(G1), .I1(P2), .Z(w44));   //: @(300,539) /sn:0 /delay:" 3" /w:[ 7 27 1 ]
  //: joint g24 (P0) @(236, 367) /w:[ 4 -1 6 3 ]
  and g39 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w15));   //: @(309,634) /sn:0 /delay:" 3" /w:[ 15 7 9 13 0 ]
  //: input g1 (Cin) @(165,285) /sn:0 /w:[ 7 ]
  //: joint g60 (G0) @(209, 627) /w:[ 14 13 -1 16 ]
  //: joint g29 (P2) @(225, 477) /w:[ 22 -1 24 21 ]
  or g51 (.I0(w42), .I1(w15), .I2(G3), .I3(w40), .I4(w39), .Z(C4));   //: @(393,655) /sn:0 /delay:" 3" /w:[ 1 1 0 1 1 1 ]
  //: joint g70 (P3) @(258, 826) /w:[ 26 25 -1 28 ]
  and g18 (.I0(P1), .I1(G0), .Z(w3));   //: @(297,411) /sn:0 /delay:" 3" /w:[ 23 7 0 ]
  //: joint g65 (G1) @(202, 668) /w:[ 10 9 -1 12 ]
  //: joint g25 (P1) @(216, 408) /w:[ 22 24 -1 21 ]
  or g10 (.I0(w2), .I1(G0), .Z(C1));   //: @(345,259) /sn:0 /delay:" 3" /w:[ 1 0 0 ]
  and g64 (.I0(G1), .I1(P2), .I2(P3), .Z(w8));   //: @(311,821) /sn:0 /delay:" 3" /w:[ 13 33 27 1 ]
  //: joint g72 (G3) @(222, 655) /w:[ 1 -1 2 4 ]
  //: joint g49 (G2) @(265, 516) /w:[ 4 -1 6 3 ]
  //: joint g50 (P3) @(258, 678) /w:[ 8 10 -1 7 ]
  //: input g6 (G2) @(165,516) /sn:0 /w:[ 7 ]
  and g68 (.I0(G2), .I1(P3), .Z(w6));   //: @(310,854) /sn:0 /delay:" 3" /w:[ 9 29 0 ]
  //: joint g58 (P3) @(258, 708) /w:[ 4 6 -1 3 ]
  //: joint g56 (P1) @(243, 632) /w:[ 6 8 -1 5 ]
  //: joint g35 (Cin) @(230, 462) /w:[ 10 9 -1 12 ]
  and g9 (.I0(P0), .I1(Cin), .Z(w2));   //: @(246,256) /sn:0 /delay:" 3" /w:[ 9 5 0 ]
  //: input g7 (P2) @(166,477) /sn:0 /w:[ 25 ]
  and g73 (.I0(P0), .I1(P1), .I2(P3), .I3(P2), .Z(PG));   //: @(310,742) /sn:0 /delay:" 3" /w:[ 17 3 0 0 0 ]
  or g71 (.I0(w4), .I1(G3), .I2(w8), .I3(w6), .Z(GG));   //: @(388,807) /sn:0 /delay:" 3" /w:[ 1 5 0 1 1 ]
  and g59 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w4));   //: @(311,784) /sn:0 /delay:" 3" /w:[ 17 0 31 23 0 ]
  //: joint g31 (G1) @(202, 385) /w:[ 2 -1 1 4 ]
  and g22 (.I0(Cin), .I1(P0), .I2(P1), .I3(P2), .Z(w45));   //: @(298,469) /sn:0 /delay:" 3" /w:[ 11 0 19 23 0 ]
  //: joint g67 (P3) @(258, 792) /w:[ 22 21 -1 24 ]
  //: joint g45 (G1) @(202, 513) /w:[ 6 5 -1 8 ]
  //: joint g41 (P1) @(243, 588) /w:[ 10 12 -1 9 ]
  //: joint g36 (P0) @(236, 467) /w:[ 1 2 -1 12 ]
  or g33 (.I0(w45), .I1(w18), .I2(w44), .I3(G2), .Z(C3));   //: @(373,508) /sn:0 /delay:" 3" /w:[ 1 1 0 5 1 ]
  //: joint g54 (P0) @(236, 583) /w:[ 14 13 -1 16 ]
  //: joint g69 (G2) @(265, 703) /w:[ 1 2 -1 8 ]
  //: output g52 (PG) @(361,742) /sn:0 /w:[ 1 ]
  //: joint g42 (P2) @(250, 593) /w:[ 12 14 -1 11 ]
  //: joint g40 (G0) @(209, 499) /w:[ 10 9 -1 12 ]
  //: joint g66 (P2) @(273, 787) /w:[ 30 29 -1 32 ]
  //: output g12 (C2) @(398,385) /sn:0 /w:[ 0 ]
  //: joint g57 (P2) @(273, 673) /w:[ 4 -1 6 3 ]
  //: joint g46 (P2) @(250, 637) /w:[ 8 10 -1 7 ]
  //: joint g28 (P1) @(216, 472) /w:[ 18 20 -1 17 ]
  and g34 (.I0(Cin), .I1(P0), .I2(P1), .I3(P2), .I4(P3), .Z(w42));   //: @(309,588) /sn:0 /anc:1 /delay:" 3" /w:[ 13 15 11 13 17 0 ]
  //: output g14 (C4) @(435,655) /sn:0 /w:[ 0 ]
  //: output g11 (C1) @(396,259) /sn:0 /w:[ 1 ]
  //: input g5 (P3) @(165,598) /sn:0 /w:[ 19 ]
  //: joint g19 (P1) @(216, 372) /w:[ 26 -1 28 25 ]
  or g21 (.I0(D8), .I1(G1), .I2(w3), .Z(C2));   //: @(359,385) /sn:0 /delay:" 3" /w:[ 1 3 1 1 ]
  //: joint g61 (P3) @(258, 745) /w:[ 1 2 -1 20 ]
  //: joint g32 (P1) @(216, 504) /w:[ 14 16 -1 13 ]
  //: joint g20 (G0) @(209, 294) /w:[ 1 -1 2 4 ]
  //: joint g43 (P3) @(258, 598) /w:[ 16 -1 18 15 ]
  //: joint g38 (P2) @(250, 509) /w:[ 16 -1 18 15 ]
  and g15 (.I0(Cin), .I1(P0), .I2(P1), .Z(D8));   //: @(298,367) /sn:0 /delay:" 3" /w:[ 0 5 27 0 ]
  //: input g0 (P0) @(164,234) /sn:0 /w:[ 11 ]
  //: joint g27 (G0) @(209, 413) /w:[ 6 5 -1 8 ]
  and g48 (.I0(G2), .I1(P3), .Z(w39));   //: @(308,706) /sn:0 /delay:" 3" /w:[ 0 5 0 ]
  //: joint g37 (P2) @(225, 509) /w:[ 19 20 -1 26 ]
  //: joint g62 (P2) @(273, 750) /w:[ 1 2 -1 28 ]
  //: joint g55 (P1) @(243, 740) /w:[ 2 4 -1 1 ]
  //: output g53 (GG) @(424,807) /sn:0 /w:[ 0 ]
  //: output g13 (C3) @(405,508) /sn:0 /w:[ 0 ]

endmodule

module signextend(Out, In);
//: interface  /sz:(183, 170) /bd:[ Li0>In[15:0](65/170) Ro0<Out[31:0](75/170) ]
input [15:0] In;    //: /sn:0 {0}(230,211)(347,211)(347,210)(463,210){1}
//: {2}(464,210)(473,210)(473,302)(614,302){3}
output [31:0] Out;    //: /sn:0 {0}(721,211)(700,211)(700,222)(620,222){1}
wire w3;    //: /sn:0 {0}(614,282)(591,282){1}
//: {2}(587,282)(572,282)(572,264){3}
//: {4}(574,262)(591,262){5}
//: {6}(595,262)(614,262){7}
//: {8}(593,264)(593,272)(614,272){9}
//: {10}(570,262)(538,262)(538,234){11}
//: {12}(540,232)(567,232){13}
//: {14}(571,232)(587,232){15}
//: {16}(591,232)(614,232){17}
//: {18}(589,234)(589,242)(614,242){19}
//: {20}(569,234)(569,252)(614,252){21}
//: {22}(536,232)(529,232)(529,120)(518,120)(518,130){23}
//: {24}(520,132)(532,132){25}
//: {26}(536,132)(542,132)(542,142)(552,142){27}
//: {28}(556,142)(567,142){29}
//: {30}(571,142)(581,142){31}
//: {32}(585,142)(614,142){33}
//: {34}(583,140)(583,130)(598,130)(598,162)(614,162){35}
//: {36}(583,144)(583,152)(614,152){37}
//: {38}(569,144)(569,172)(614,172){39}
//: {40}(554,140)(554,130)(577,130)(577,192)(614,192){41}
//: {42}(554,144)(554,182)(614,182){43}
//: {44}(534,130)(534,120)(549,120)(549,212)(614,212){45}
//: {46}(534,134)(534,202)(614,202){47}
//: {48}(516,132)(464,132)(464,205){49}
//: {50}(518,134)(518,222)(614,222){51}
//: {52}(589,284)(589,292)(614,292){53}
//: enddecls

  //: joint g8 (w3) @(589, 232) /w:[ 16 -1 15 18 ]
  //: joint g4 (w3) @(569, 142) /w:[ 30 -1 29 38 ]
  //: joint g3 (w3) @(583, 142) /w:[ 32 34 31 36 ]
  tran g2(.Z(w3), .I(In[15]));   //: @(464,208) /sn:0 /R:1 /w:[ 49 1 2 ] /ss:0
  concat g1 (.I0(In), .I1(w3), .I2(w3), .I3(w3), .I4(w3), .I5(w3), .I6(w3), .I7(w3), .I8(w3), .I9(w3), .I10(w3), .I11(w3), .I12(w3), .I13(w3), .I14(w3), .I15(w3), .I16(w3), .Z(Out));   //: @(619,222) /sn:0 /w:[ 3 53 0 9 7 21 19 17 51 45 47 41 43 39 35 37 33 1 ] /dr:0
  //: joint g10 (w3) @(538, 232) /w:[ 12 -1 22 11 ]
  //: joint g6 (w3) @(534, 132) /w:[ 26 44 25 46 ]
  //: joint g9 (w3) @(569, 232) /w:[ 14 -1 13 20 ]
  //: joint g7 (w3) @(518, 132) /w:[ 24 23 48 50 ]
  //: joint g12 (w3) @(572, 262) /w:[ 4 -1 10 3 ]
  //: output g14 (Out) @(718,211) /sn:0 /w:[ 0 ]
  //: joint g11 (w3) @(593, 262) /w:[ 6 -1 5 8 ]
  //: joint g5 (w3) @(554, 142) /w:[ 28 40 27 42 ]
  //: input g0 (In) @(228,211) /sn:0 /w:[ 0 ]
  //: joint g13 (w3) @(589, 282) /w:[ 1 -1 2 52 ]

endmodule

module fetch(reset, clk, Inst, PCNext, PCNew);
//: interface  /sz:(420, 354) /bd:[ Li0>PCNew[31:0](181/354) Li1>reset(96/354) Li2>clk(262/354) Ro0<Inst[31:0](271/354) Ro1<PCNext[31:0](49/354) ]
supply0 w4;    //: /sn:0 {0}(258,62)(258,93)(257,93)(257,101){1}
input [31:0] PCNew;    //: /sn:0 {0}(241,139)(231,139)(231,138)(163,138){1}
output [31:0] Inst;    //: /sn:0 /dp:1 {0}(366,149)(468,149)(468,137)(574,137){1}
output [31:0] PCNext;    //: /sn:0 /dp:1 {0}(436,68)(541,68)(541,65)(551,65){1}
supply0 w1;    //: /sn:0 {0}(353,202)(353,195)(349,195)(349,176){1}
input clk;    //: /sn:0 {0}(61,183)(196,183)(196,189)(252,189)(252,177){1}
supply0 w2;    //: /sn:0 {0}(419,-6)(419,37)(421,37)(421,44){1}
input reset;    //: /sn:0 {0}(151,75)(189,75){1}
//: {2}(193,75)(247,75)(247,101){3}
//: {4}(191,73)(191,63)(194,63)(194,33){5}
wire w7;    //: /sn:0 {0}(421,92)(421,121){1}
wire [31:0] w0;    //: /sn:0 {0}(262,139)(289,139){1}
//: {2}(293,139)(310,139)(310,151)(331,151){3}
//: {4}(291,137)(291,52)(407,52){5}
wire [31:0] w3;    //: /sn:0 {0}(382,80)(397,80)(397,84)(407,84){1}
//: enddecls

  add g8 (.A(w3), .B(w0), .S(PCNext), .CI(w2), .CO(w7));   //: @(423,68) /sn:0 /R:1 /w:[ 1 5 0 1 0 ]
  led g4 (.I(reset));   //: @(194,26) /sn:0 /w:[ 5 ] /type:0
  register g3 (.Q(w0), .D(PCNew), .EN(w4), .CLR(!reset), .CK(!clk));   //: @(252,139) /sn:0 /R:1 /w:[ 0 0 1 3 1 ]
  //: input g2 (reset) @(149,75) /sn:0 /w:[ 0 ]
  //: input g1 (clk) @(59,183) /sn:0 /w:[ 0 ]
  //: dip g10 (w3) @(344,80) /sn:0 /R:1 /w:[ 0 ] /st:1
  //: output g6 (Inst) @(571,137) /sn:0 /w:[ 1 ]
  //: supply0 g7 (w4) @(258,56) /sn:0 /R:2 /w:[ 0 ]
  //: joint g9 (w0) @(291, 139) /w:[ 2 4 1 -1 ]
  //: supply0 g12 (w2) @(419,-12) /sn:0 /R:2 /w:[ 0 ]
  //: supply0 g5 (w1) @(353,208) /sn:0 /w:[ 0 ]
  //: output g11 (PCNext) @(548,65) /sn:0 /w:[ 1 ]
  //: joint g14 (reset) @(191, 75) /w:[ 2 4 1 -1 ]
  //: input g0 (PCNew) @(161,138) /sn:0 /w:[ 1 ]
  rom g13 (.A(w0), .D(Inst), .OE(w1));   //: @(349,150) /w:[ 3 0 1 ]

endmodule

module CLA16Bits(B, Cin, A, GG, Cout, PG, S);
//: interface  /sz:(322, 143) /bd:[ Ti0>A[15:0](70/322) Ti1>B[15:0](209/322) Ri0>Cin(75/143) Lo0<PG(111/143) Lo1<GG(58/143) Bo0<Cout[15:0](182/322) Bo1<S[15:0](235/322) ]
input [15:0] B;    //: /sn:0 {0}(-203,-33)(-70,-33){1}
//: {2}(-69,-33)(191,-33){3}
//: {4}(192,-33)(463,-33){5}
//: {6}(464,-33)(723,-33){7}
//: {8}(724,-33)(877,-33){9}
output GG;    //: /sn:0 /dp:1 {0}(693,354)(693,421){1}
input [15:0] A;    //: /sn:0 {0}(875,-108)(686,-108){1}
//: {2}(685,-108)(415,-108){3}
//: {4}(414,-108)(157,-108){5}
//: {6}(156,-108)(-107,-108){7}
//: {8}(-108,-108)(-201,-108){9}
output PG;    //: /sn:0 /dp:1 {0}(541,354)(541,419){1}
input Cin;    //: /sn:0 {0}(826,93)(971,93)(971,94){1}
//: {2}(973,96)(979,96)(979,87)(989,87){3}
//: {4}(971,98)(971,324)(831,324){5}
output Cout;    //: /sn:0 /dp:1 {0}(-145,312)(-265,312)(-265,316)(-255,316){1}
output [15:0] S;    //: /sn:0 /dp:1 {0}(885,194)(925,194){1}
wire w16;    //: /sn:0 {0}(802,266)(802,232)(750,232)(750,156){1}
wire w6;    //: /sn:0 {0}(294,90)(361,90)(361,266){1}
wire [3:0] w7;    //: /sn:0 {0}(155,153)(155,189)(879,189){1}
wire w25;    //: /sn:0 /dp:1 {0}(98,266)(98,82)(32,82){1}
wire [3:0] w39;    //: /sn:0 {0}(687,156)(687,209)(879,209){1}
wire w22;    //: /sn:0 {0}(38,266)(38,223)(-44,223)(-44,145){1}
wire [3:0] w0;    //: /sn:0 /dp:1 {0}(157,-104)(157,-83)(155,-83)(155,55){1}
wire [3:0] w36;    //: /sn:0 {0}(687,58)(687,46)(686,46)(686,-104){1}
wire w20;    //: /sn:0 {0}(313,266)(313,234)(218,234)(218,153){1}
wire [3:0] w37;    //: /sn:0 {0}(724,58)(724,-29){1}
wire w18;    //: /sn:0 {0}(566,266)(566,252)(486,252)(486,157){1}
wire w19;    //: /sn:0 {0}(513,266)(513,167)(529,167)(529,157){1}
wire w12;    //: /sn:0 {0}(562,94)(602,94)(602,266){1}
wire w23;    //: /sn:0 {0}(-24,266)(-24,250)(-1,250)(-1,145){1}
wire [3:0] w10;    //: /sn:0 {0}(423,59)(423,33)(415,33)(415,-104){1}
wire [3:0] w1;    //: /sn:0 /dp:1 {0}(192,-29)(192,55){1}
wire [3:0] w31;    //: /sn:0 /dp:1 {0}(879,199)(423,199)(423,157){1}
wire w17;    //: /sn:0 {0}(743,266)(743,241)(791,241)(791,156){1}
wire [3:0] w27;    //: /sn:0 /dp:1 {0}(464,-29)(464,49)(460,49)(460,59){1}
wire [3:0] w14;    //: /sn:0 /dp:1 {0}(-107,-104)(-107,47){1}
wire [3:0] w2;    //: /sn:0 {0}(-70,47)(-70,-21)(-69,-21)(-69,-29){1}
wire [3:0] w26;    //: /sn:0 /dp:1 {0}(879,179)(-107,179)(-107,145){1}
wire w9;    //: /sn:0 /dp:1 {0}(261,153)(261,256)(258,256)(258,266){1}
//: enddecls

  CLL g4 (.P3(w23), .G3(w22), .P2(w9), .G2(w20), .P1(w19), .G1(w18), .P0(w17), .G0(w16), .Cin(Cin), .C3(w25), .C2(w6), .C1(w12), .C4(Cout), .PG(PG), .GG(GG));   //: @(-144, 267) /sz:(974, 86) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>5 To0<0 To1<1 To2<1 Lo0<0 Bo0<0 Bo1<0 ]
  tran g8(.Z(w36), .I(A[3:0]));   //: @(686,-110) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g16(.Z(w14), .I(A[15:12]));   //: @(-107,-110) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  CLA g3 (.B(w37), .A(w36), .Cin(Cin), .p0(w17), .g0(w16), .S(w39));   //: @(663, 59) /sz:(162, 96) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Bo0<1 Bo1<1 Bo2<0 ]
  tran g17(.Z(w1), .I(B[11:8]));   //: @(192,-35) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  CLA g2 (.B(w27), .A(w10), .Cin(w12), .p0(w19), .g0(w18), .S(w31));   //: @(399, 60) /sz:(162, 96) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>0 Bo0<1 Bo1<1 Bo2<1 ]
  CLA g1 (.B(w1), .A(w0), .Cin(w6), .p0(w9), .g0(w20), .S(w7));   //: @(131, 56) /sz:(162, 96) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<0 Bo1<1 Bo2<0 ]
  tran g18(.Z(w27), .I(B[7:4]));   //: @(464,-35) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g10(.Z(w0), .I(A[11:8]));   //: @(157,-110) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  //: input g6 (B) @(-205,-33) /sn:0 /w:[ 0 ]
  tran g7(.Z(w37), .I(B[3:0]));   //: @(724,-35) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g9(.Z(w10), .I(A[7:4]));   //: @(415,-110) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  concat g12 (.I0(w39), .I1(w31), .I2(w7), .I3(w26), .Z(S));   //: @(884,194) /sn:0 /w:[ 1 0 1 0 0 ] /dr:0
  //: input g14 (Cin) @(991,87) /sn:0 /R:2 /w:[ 3 ]
  //: input g5 (A) @(-203,-108) /sn:0 /w:[ 9 ]
  tran g11(.Z(w2), .I(B[15:12]));   //: @(-69,-35) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: output g19 (GG) @(693,418) /sn:0 /R:3 /w:[ 1 ]
  //: output g21 (Cout) @(-258,316) /sn:0 /w:[ 1 ]
  //: output g20 (PG) @(541,416) /sn:0 /R:3 /w:[ 1 ]
  CLA g0 (.B(w2), .A(w14), .Cin(w25), .p0(w23), .g0(w22), .S(w26));   //: @(-131, 48) /sz:(162, 96) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>1 Bo0<1 Bo1<1 Bo2<1 ]
  //: joint g15 (Cin) @(971, 96) /w:[ 2 1 -1 4 ]
  //: output g13 (S) @(922,194) /sn:0 /w:[ 1 ]

endmodule

module PFA(Pi, S, Ci, B, Gi, A);
//: interface  /sz:(77, 43) /bd:[ Ti0>A(15/77) Ti1>B(44/77) Ti2>Ci(71/77) Ti3>A(14/77) Ti4>B(43/77) Ti5>Ci(70/77) Ti6>APFA(13/77) Ti7>BPFA(62/77) Ri0>CinPFA(20/43) Bo0<S(23/77) Bo1<Pi(50/77) Bo2<Gi(71/77) Bo3<S(22/77) Bo4<Pi(49/77) Bo5<Gi(70/77) Bo6<PPFA(8/77) Bo7<GFPA(20/77) Bo8<SPFA(65/77) ]
input B;    //: /sn:0 {0}(206,145)(223,145){1}
//: {2}(227,145)(269,145)(269,133)(279,133){3}
//: {4}(225,147)(225,188){5}
//: {6}(227,190)(354,190){7}
//: {8}(225,192)(225,229)(356,229){9}
output Gi;    //: /sn:0 {0}(435,225)(387,225)(387,227)(377,227){1}
input A;    //: /sn:0 {0}(205,117)(246,117){1}
//: {2}(250,117)(269,117)(269,128)(279,128){3}
//: {4}(248,119)(248,183){5}
//: {6}(250,185)(354,185){7}
//: {8}(248,187)(248,224)(356,224){9}
output Pi;    //: /sn:0 /dp:1 {0}(375,188)(422,188)(422,187)(432,187){1}
input Ci;    //: /sn:0 /dp:1 {0}(352,146)(315,146)(315,174)(204,174){1}
output S;    //: /sn:0 /dp:1 {0}(373,144)(424,144)(424,145)(433,145){1}
wire w2;    //: /sn:0 {0}(300,131)(342,131)(342,141)(352,141){1}
//: enddecls

  //: output g4 (Pi) @(429,187) /sn:0 /w:[ 1 ]
  or g8 (.I0(A), .I1(B), .Z(Pi));   //: @(365,188) /sn:0 /delay:" 3" /w:[ 7 7 0 ]
  //: output g3 (S) @(430,145) /sn:0 /w:[ 1 ]
  //: input g2 (Ci) @(202,174) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(204,145) /sn:0 /w:[ 0 ]
  //: joint g10 (A) @(248, 117) /w:[ 2 -1 1 4 ]
  xor g6 (.I0(A), .I1(B), .Z(w2));   //: @(290,131) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  xor g7 (.I0(w2), .I1(Ci), .Z(S));   //: @(363,144) /sn:0 /delay:" 4" /w:[ 1 0 0 ]
  and g9 (.I0(A), .I1(B), .Z(Gi));   //: @(367,227) /sn:0 /delay:" 3" /w:[ 9 9 1 ]
  //: joint g12 (B) @(225, 145) /w:[ 2 -1 1 4 ]
  //: output g5 (Gi) @(432,225) /sn:0 /w:[ 0 ]
  //: joint g11 (A) @(248, 185) /w:[ 6 5 -1 8 ]
  //: input g0 (A) @(203,117) /sn:0 /w:[ 0 ]
  //: joint g13 (B) @(225, 190) /w:[ 6 5 -1 8 ]

endmodule

module CSA16bits(Cin, B, S, A, Cout);
//: interface  /sz:(257, 128) /bd:[ Ti0>A[15:0](61/257) Ti1>B[15:0](178/257) Ri0>Cin(70/128) Bo0<S[15:0](165/257) Bo1<Cout(52/257) ]
input [15:0] B;    //: /sn:0 {0}(961,126)(834,126){1}
//: {2}(833,126)(748,126){3}
//: {4}(747,126)(670,126){5}
//: {6}(669,126)(585,126){7}
//: {8}(584,126)(429,126){9}
//: {10}(428,126)(247,126){11}
//: {12}(246,126)(80,126){13}
//: {14}(79,126)(-26,126){15}
input [15:0] A;    //: /sn:0 {0}(-25,166)(58,166){1}
//: {2}(59,166)(224,166){3}
//: {4}(225,166)(403,166){5}
//: {6}(404,166)(601,166){7}
//: {8}(602,166)(685,166){9}
//: {10}(686,166)(762,166){11}
//: {12}(763,166)(849,166){13}
//: {14}(850,166)(962,166){15}
input Cin;    //: /sn:0 {0}(917,269)(865,269){1}
output Cout;    //: /sn:0 /dp:1 {0}(146,235)(146,221)(11,221){1}
output [15:0] S;    //: /sn:0 /dp:1 {0}(885,432)(1019,432)(1019,404)(1029,404){1}
wire w16;    //: /sn:0 {0}(585,246)(585,130){1}
wire [3:0] w6;    //: /sn:0 {0}(247,236)(247,130){1}
wire w7;    //: /sn:0 {0}(291,236)(291,205)(504,205)(504,235){1}
wire w34;    //: /sn:0 {0}(849,291)(849,507)(879,507){1}
wire w25;    //: /sn:0 {0}(778,267)(788,267)(788,304)(832,304)(832,291){1}
wire [3:0] w4;    //: /sn:0 {0}(98,235)(98,217)(115,217)(115,234)(108,234)(108,312)(96,312)(96,335){1}
//: {2}(96,336)(96,350){3}
//: {4}(96,351)(96,359)(95,359)(95,367){5}
//: {6}(95,368)(95,378)(94,378)(94,388){7}
//: {8}(94,389)(94,394){9}
wire w3;    //: /sn:0 {0}(299,374)(299,380){1}
//: {2}(297,382)(280,382)(280,381)(272,381){3}
//: {4}(299,384)(299,397)(879,397){5}
wire w36;    //: /sn:0 {0}(879,427)(273,427){1}
wire w22;    //: /sn:0 {0}(686,247)(686,170){1}
wire [3:0] w0;    //: /sn:0 {0}(59,235)(59,170){1}
wire w20;    //: /sn:0 {0}(700,267)(710,267)(710,299)(745,299)(745,289){1}
wire w30;    //: /sn:0 {0}(879,457)(475,457)(475,445)(467,445){1}
wire w42;    //: /sn:0 {0}(879,367)(126,367)(126,356){1}
//: {2}(126,352)(126,347){3}
//: {4}(124,354)(108,354)(108,351)(100,351){5}
wire w37;    //: /sn:0 {0}(879,417)(280,417)(280,410)(272,410){1}
wire w18;    //: /sn:0 {0}(879,487)(684,487)(684,289){1}
wire w19;    //: /sn:0 {0}(599,288)(599,477)(879,477){1}
wire w12;    //: /sn:0 {0}(483,235)(483,218)(549,218)(549,298)(582,298)(582,288){1}
wire [3:0] w10;    //: /sn:0 {0}(404,235)(404,170){1}
wire w21;    //: /sn:0 {0}(670,247)(670,130){1}
wire w31;    //: /sn:0 {0}(835,249)(835,138)(834,138)(834,130){1}
wire [3:0] w1;    //: /sn:0 {0}(80,235)(80,130){1}
wire w32;    //: /sn:0 {0}(851,249)(851,178)(850,178)(850,170){1}
wire w8;    //: /sn:0 /dp:1 {0}(879,497)(762,497)(762,289){1}
wire w17;    //: /sn:0 {0}(601,246)(601,178)(602,178)(602,170){1}
wire w27;    //: /sn:0 {0}(764,247)(764,178)(763,178)(763,170){1}
wire w35;    //: /sn:0 {0}(879,437)(573,437)(573,383){1}
//: {2}(573,379)(573,365){3}
//: {4}(571,381)(457,381)(457,383)(453,383){5}
wire w33;    //: /sn:0 {0}(494,436)(493,436){1}
//: {2}(491,434)(491,421)(453,421){3}
//: {4}(491,438)(491,447)(879,447){5}
wire w28;    //: /sn:0 {0}(879,467)(475,467)(475,465)(467,465){1}
wire [3:0] w14;    //: /sn:0 {0}(456,235)(456,217)(442,217)(442,341)(449,341)(449,382){1}
//: {2}(449,383)(449,420){3}
//: {4}(449,421)(449,431)(463,431)(463,444){5}
//: {6}(463,445)(463,464){7}
//: {8}(463,465)(463,472){9}
wire w41;    //: /sn:0 {0}(879,377)(107,377)(107,368)(99,368){1}
wire w2;    //: /sn:0 {0}(124,235)(124,217)(313,217)(313,236){1}
wire [3:0] w11;    //: /sn:0 {0}(428,235)(428,138)(429,138)(429,130){1}
wire w15;    //: /sn:0 {0}(615,266)(630,266)(630,299)(667,299)(667,289){1}
wire w38;    //: /sn:0 {0}(879,407)(287,407)(287,397){1}
//: {2}(287,393)(287,391){3}
//: {4}(285,395)(272,395){5}
wire [3:0] w5;    //: /sn:0 {0}(226,236)(226,178)(225,178)(225,170){1}
wire w43;    //: /sn:0 {0}(879,357)(146,357)(146,343){1}
//: {2}(146,339)(146,337){3}
//: {4}(144,341)(108,341)(108,336)(100,336){5}
wire w26;    //: /sn:0 {0}(748,247)(748,130){1}
wire [3:0] w9;    //: /sn:0 {0}(265,236)(265,218)(279,218)(279,334)(268,334)(268,380){1}
//: {2}(268,381)(268,394){3}
//: {4}(268,395)(268,409){5}
//: {6}(268,410)(268,418)(269,418)(269,426){7}
//: {8}(269,427)(269,436){9}
wire w40;    //: /sn:0 {0}(879,387)(106,387)(106,389)(98,389){1}
//: enddecls

  tran g44(.Z(w43), .I(w4[3]));   //: @(94,336) /sn:0 /R:2 /w:[ 5 2 1 ] /ss:1
  //: input g8 (Cin) @(919,269) /sn:0 /R:2 /w:[ 0 ]
  FA g4 (.A(w22), .B(w21), .Cin(w20), .S(w18), .Cout(w15));   //: @(659, 248) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Bo0<1 Bo1<1 ]
  tran g16(.Z(w0), .I(A[15:12]));   //: @(59,164) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  FA g3 (.A(w17), .B(w16), .Cin(w15), .S(w19), .Cout(w12));   //: @(574, 247) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Bo0<0 Bo1<1 ]
  tran g26(.Z(w28), .I(w14[0]));   //: @(461,465) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  //: input g17 (B) @(963,126) /sn:0 /R:2 /w:[ 0 ]
  CSA g2 (.Cin(w12), .B(w11), .A(w10), .S(w14), .Cout(w7));   //: @(395, 236) /sz:(127, 64) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 To0<0 To1<1 ]
  //: joint g30 (w35) @(573, 381) /w:[ -1 2 4 1 ]
  tran g23(.Z(w6), .I(B[11:8]));   //: @(247,124) /sn:0 /R:1 /w:[ 1 12 11 ] /ss:1
  tran g39(.Z(w40), .I(w4[0]));   //: @(92,389) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  tran g24(.Z(w1), .I(B[15:12]));   //: @(80,124) /sn:0 /R:1 /w:[ 1 14 13 ] /ss:1
  CSA g1 (.Cin(w7), .B(w6), .A(w5), .S(w9), .Cout(w2));   //: @(217, 237) /sz:(127, 64) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 To0<0 To1<1 ]
  tran g29(.Z(w33), .I(w14[2]));   //: @(447,421) /sn:0 /R:2 /w:[ 3 4 3 ] /ss:1
  tran g18(.Z(w31), .I(B[0]));   //: @(834,124) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  //: output g25 (S) @(1026,404) /sn:0 /w:[ 1 ]
  tran g10(.Z(w32), .I(A[0]));   //: @(850,164) /sn:0 /R:1 /w:[ 1 13 14 ] /ss:1
  FA g6 (.A(w32), .B(w31), .Cin(Cin), .S(w34), .Cout(w25));   //: @(824, 250) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<1 ]
  //: joint g35 (w38) @(287, 395) /w:[ -1 2 4 1 ]
  //: input g9 (A) @(964,166) /sn:0 /R:2 /w:[ 15 ]
  //: output g7 (Cout) @(14,221) /sn:0 /R:2 /w:[ 1 ]
  tran g31(.Z(w35), .I(w14[3]));   //: @(447,383) /sn:0 /R:2 /w:[ 5 2 1 ] /ss:1
  tran g22(.Z(w11), .I(B[7:4]));   //: @(429,124) /sn:0 /R:1 /w:[ 1 10 9 ] /ss:1
  //: joint g41 (w42) @(126, 354) /w:[ -1 2 4 1 ]
  tran g36(.Z(w38), .I(w9[2]));   //: @(266,395) /sn:0 /R:2 /w:[ 5 4 3 ] /ss:1
  concat g33 (.I0(w34), .I1(w8), .I2(w18), .I3(w19), .I4(w28), .I5(w30), .I6(w33), .I7(w35), .I8(w36), .I9(w37), .I10(w38), .I11(w3), .I12(w40), .I13(w41), .I14(w42), .I15(w43), .Z(S));   //: @(884,432) /sn:0 /w:[ 1 0 0 1 0 0 5 0 0 0 0 5 0 0 0 0 0 ] /dr:0
  tran g42(.Z(w42), .I(w4[2]));   //: @(94,351) /sn:0 /R:2 /w:[ 5 4 3 ] /ss:1
  tran g40(.Z(w41), .I(w4[1]));   //: @(93,368) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1
  tran g12(.Z(w22), .I(A[2]));   //: @(686,164) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:1
  tran g34(.Z(w37), .I(w9[1]));   //: @(266,410) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1
  //: joint g28 (w33) @(491, 436) /w:[ 1 2 -1 4 ]
  tran g14(.Z(w10), .I(A[7:4]));   //: @(404,164) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g11(.Z(w27), .I(A[1]));   //: @(763,164) /sn:0 /R:1 /w:[ 1 11 12 ] /ss:1
  FA g5 (.A(w27), .B(w26), .Cin(w25), .S(w8), .Cout(w20));   //: @(737, 248) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Bo0<1 Bo1<1 ]
  tran g21(.Z(w16), .I(B[3]));   //: @(585,124) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  tran g19(.Z(w26), .I(B[1]));   //: @(748,124) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g32(.Z(w36), .I(w9[0]));   //: @(267,427) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  tran g20(.Z(w21), .I(B[2]));   //: @(670,124) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  //: joint g43 (w43) @(146, 341) /w:[ -1 2 4 1 ]
  tran g38(.Z(w3), .I(w9[3]));   //: @(266,381) /sn:0 /R:2 /w:[ 3 2 1 ] /ss:1
  tran g15(.Z(w5), .I(A[11:8]));   //: @(225,164) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  CSA g0 (.Cin(w2), .B(w1), .A(w0), .S(w4), .Cout(Cout));   //: @(50, 236) /sz:(127, 64) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 To0<0 To1<0 ]
  tran g27(.Z(w30), .I(w14[1]));   //: @(461,445) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1
  //: joint g37 (w3) @(299, 382) /w:[ -1 1 2 4 ]
  tran g13(.Z(w17), .I(A[3]));   //: @(602,164) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1

endmodule

module Regs8x324(SB, SA, BOUT, AOUT, Pop, clr, clk, RegWr, SD, DIN);
//: interface  /sz:(98, 69) /bd:[ Ti0>DIN[31:0](47/98) Ti1>Pop(85/98) Ti2>DIN[31:0](47/98) Li0>SD[2:0](35/69) Li1>SA[2:0](11/69) Li2>SB[2:0](22/69) Li3>RegWr(47/69) Li4>clk(59/69) Li5>SD[2:0](35/69) Li6>SA[2:0](11/69) Li7>SB[2:0](22/69) Li8>RegWr(47/69) Li9>clk(59/69) Ri0>clr(35/69) Ri1>clr(35/69) Bo0<AOUT[31:0](37/98) Bo1<BOUT[31:0](65/98) Bo2<AOUT[31:0](37/98) Bo3<BOUT[31:0](65/98) ]
supply0 w13;    //: /sn:0 /dp:1 {0}(947,500)(947,469){1}
input Pop;    //: /sn:0 {0}(1019,286)(949,286)(949,295){1}
//: {2}(947,297)(744,297)(744,299){3}
//: {4}(742,301)(685,301)(685,294)(659,294){5}
//: {6}(744,303)(744,426){7}
//: {8}(949,299)(949,379){9}
input [31:0] DIN;    //: /sn:0 {0}(531,269)(531,318){1}
//: {2}(533,320)(715,320){3}
//: {4}(719,320)(807,320)(807,365){5}
//: {6}(809,367)(915,367){7}
//: {8}(919,367)(969,367)(969,364)(977,364){9}
//: {10}(979,362)(979,351){11}
//: {12}(979,366)(979,392)(965,392){13}
//: {14}(917,369)(917,508)(933,508){15}
//: {16}(807,369)(807,429){17}
//: {18}(717,322)(717,352){19}
//: {20}(529,320)(435,320){21}
//: {22}(431,320)(342,320){23}
//: {24}(338,320)(264,320){25}
//: {26}(260,320)(181,320)(181,352){27}
//: {28}(262,322)(262,439){29}
//: {30}(340,322)(340,351){31}
//: {32}(433,322)(433,436){33}
//: {34}(531,322)(531,348){35}
output [31:0] BOUT;    //: /sn:0 {0}(516,697)(516,672){1}
input [2:0] SD;    //: /sn:0 {0}(782,138)(852,138)(852,156){1}
input [2:0] SB;    //: /sn:0 {0}(466,659)(493,659){1}
supply1 w21;    //: /sn:0 {0}(828,169)(801,169)(801,153){1}
input RegWr;    //: /sn:0 {0}(48,363)(68,363)(68,378)(82,378){1}
input clr;    //: /sn:0 /dp:1 {0}(959,337)(1032,337){1}
input [2:0] SA;    //: /sn:0 {0}(256,657)(231,657){1}
input clk;    //: /sn:0 {0}(82,383)(68,383)(68,398)(55,398){1}
output [31:0] AOUT;    //: /sn:0 {0}(279,670)(279,702){1}
wire [31:0] w6;    //: /sn:0 /dp:1 {0}(936,402)(629,402)(629,433){1}
wire w16;    //: /sn:0 {0}(638,296)(542,296)(542,454)(552,454){1}
wire w7;    //: /sn:0 {0}(472,451)(513,451)(513,405)(848,405)(848,185){1}
wire w4;    //: /sn:0 {0}(943,337)(906,337){1}
//: {2}(902,337)(767,337){3}
//: {4}(763,337)(588,337){5}
//: {6}(584,337)(390,337){7}
//: {8}(386,337)(231,337)(231,357)(220,357){9}
//: {10}(388,339)(388,356)(379,356){11}
//: {12}(586,339)(586,353)(570,353){13}
//: {14}(765,339)(765,357)(756,357){15}
//: {16}(904,339)(904,417)(865,417){17}
//: {18}(861,417)(675,417){19}
//: {20}(671,417)(489,417){21}
//: {22}(485,417)(302,417)(302,444)(301,444){23}
//: {24}(487,419)(487,441)(472,441){25}
//: {26}(673,419)(673,438)(668,438){27}
//: {28}(863,419)(863,434)(846,434){29}
wire w3;    //: /sn:0 {0}(835,185)(835,397)(330,397)(330,454)(301,454){1}
wire w0;    //: /sn:0 {0}(552,459)(542,459)(542,479){1}
//: {2}(544,481)(764,481)(764,439)(770,439){3}
//: {4}(540,481)(390,481){5}
//: {6}(388,479)(388,446)(396,446){7}
//: {8}(386,481)(214,481){9}
//: {10}(212,479)(212,449)(225,449){11}
//: {12}(210,481)(125,481)(125,383){13}
//: {14}(127,381)(291,381){15}
//: {16}(295,381)(477,381){17}
//: {18}(481,381)(635,381){19}
//: {20}(639,381)(662,381)(662,362)(680,362){21}
//: {22}(637,379)(637,314)(669,314)(669,299)(659,299){23}
//: {24}(479,379)(479,358)(494,358){25}
//: {26}(293,379)(293,361)(303,361){27}
//: {28}(125,379)(125,362)(144,362){29}
//: {30}(123,381)(103,381){31}
wire [31:0] R2;    //: {0}(262,641)(262,537){1}
//: {2}(264,535)(499,535)(499,643){3}
//: {4}(262,533)(262,502){5}
//: {6}(262,498)(262,460){7}
//: {8}(260,500)(68,500)(68,512)(53,512)(53,502){9}
wire [31:0] R7;    //: {0}(807,450)(807,609)(541,609){1}
//: {2}(537,609)(302,609)(302,641){3}
//: {4}(539,611)(539,643){5}
wire w20;    //: /sn:0 {0}(861,185)(861,390)(749,390)(749,426){1}
wire w12;    //: /sn:0 {0}(756,367)(787,367)(787,258)(868,258)(868,185){1}
wire w19;    //: /sn:0 /dp:1 {0}(668,448)(731,448)(731,457)(746,457)(746,447){1}
wire w10;    //: /sn:0 {0}(846,444)(875,444)(875,185){1}
wire [31:0] R4;    //: {0}(340,372)(340,545){1}
//: {2}(342,547)(505,547)(505,643){3}
//: {4}(338,547)(268,547)(268,641){5}
wire [31:0] R5a1;    //: /dp:3 {0}(288,641)(288,586)(525,586){1}
//: {2}(529,586)(629,586)(629,539){3}
//: {4}(631,537)(755,537)(755,694)(770,694)(770,684){5}
//: {6}(629,535)(629,454){7}
//: {8}(527,588)(527,617)(525,617)(525,643){9}
wire w1;    //: /sn:0 /dp:1 {0}(946,584)(946,558)(947,558)(947,548){1}
wire [31:0] R3;    //: {0}(512,643)(512,559)(435,559){1}
//: {2}(433,557)(433,457){3}
//: {4}(431,559)(275,559)(275,641){5}
wire w8;    //: /sn:0 {0}(220,367)(249,367)(249,213)(828,213)(828,185){1}
wire [31:0] R0t1;    //: /dp:3 {0}(492,643)(492,523)(257,523){1}
//: {2}(253,523)(181,523)(181,419){3}
//: {4}(181,415)(181,373){5}
//: {6}(179,417)(119,417)(119,290){7}
//: {8}(255,525)(255,641){9}
wire w14;    //: /sn:0 {0}(379,366)(414,366)(414,229)(841,229)(841,185){1}
wire [31:0] w2;    //: /sn:0 /dp:1 {0}(920,592)(927,592)(927,540)(933,540){1}
wire [31:0] R4a0;    //: /sn:0 {0}(531,369)(531,427){1}
//: {2}(533,429)(572,429)(572,190){3}
//: {4}(531,431)(531,574)(520,574){5}
//: {6}(516,574)(282,574)(282,641){7}
//: {8}(518,576)(518,587)(519,587)(519,643){9}
wire w15;    //: /sn:0 {0}(570,363)(608,363)(608,244)(855,244)(855,185){1}
wire [31:0] R10;    //: /sn:0 {0}(295,641)(295,600)(530,600){1}
//: {2}(534,600)(717,600)(717,373){3}
//: {4}(532,602)(532,643){5}
wire w5;    //: /sn:0 /dp:1 {0}(592,443)(583,443)(583,457)(573,457){1}
wire [31:0] w9;    //: /sn:0 /dp:1 {0}(962,524)(970,524)(970,412)(965,412){1}
//: enddecls

  //: input g4 (SB) @(464,659) /sn:0 /w:[ 0 ]
  //: joint g8 (R4a0) @(518, 574) /w:[ 5 -1 6 8 ]
  led g44 (.I(R4a0));   //: @(572,183) /sn:0 /w:[ 3 ] /type:2
  //: joint g16 (R3) @(433, 559) /w:[ 1 2 4 -1 ]
  //: input g3 (SA) @(229,657) /sn:0 /w:[ 1 ]
  //: dip g47 (w2) @(882,592) /sn:0 /R:1 /w:[ 0 ] /st:1
  //: joint g26 (DIN) @(340, 320) /w:[ 23 -1 24 30 ]
  //: joint g17 (R4) @(340, 547) /w:[ 2 1 4 -1 ]
  //: output g2 (BOUT) @(516,694) /sn:0 /R:3 /w:[ 0 ]
  register R5 (.Q(R5a1), .D(w6), .EN(w19), .CLR(w4), .CK(!w5));   //: @(629,443) /w:[ 7 1 0 27 0 ]
  //: joint g30 (w0) @(212, 481) /w:[ 9 10 12 -1 ]
  //: joint g23 (w4) @(765, 337) /w:[ 3 -1 4 14 ]
  //: joint g24 (DIN) @(531, 320) /w:[ 2 1 20 34 ]
  //: joint g39 (DIN) @(262, 320) /w:[ 25 -1 26 28 ]
  //: output g1 (AOUT) @(279,699) /sn:0 /R:3 /w:[ 1 ]
  //: joint g29 (w0) @(388, 481) /w:[ 5 6 8 -1 ]
  or g60 (.I0(w16), .I1(w0), .Z(w5));   //: @(563,457) /sn:0 /w:[ 1 0 1 ]
  register R2 (.Q(R4), .D(DIN), .EN(w14), .CLR(w4), .CK(!w0));   //: @(340,361) /w:[ 0 31 0 11 27 ]
  //: joint g51 (DIN) @(979, 364) /w:[ -1 10 9 12 ]
  //: joint g18 (R2) @(262, 535) /w:[ 2 4 -1 1 ]
  register R7 (.Q(R7), .D(DIN), .EN(w10), .CLR(w4), .CK(!w0));   //: @(807,439) /w:[ 0 17 0 29 3 ]
  not g25 (.I(clr), .Z(w4));   //: @(953,337) /sn:0 /R:2 /w:[ 0 0 ]
  //: supply1 g10 (w21) @(812,153) /sn:0 /w:[ 1 ]
  //: input g49 (Pop) @(1021,286) /sn:0 /R:2 /w:[ 0 ]
  register R6 (.Q(R10), .D(DIN), .EN(w12), .CLR(w4), .CK(!w0));   //: @(717,362) /w:[ 3 19 0 15 21 ]
  //: joint g6 (R7) @(539, 609) /w:[ 1 -1 2 4 ]
  mux g50 (.I0(DIN), .I1(w9), .S(Pop), .Z(w6));   //: @(949,402) /sn:0 /R:3 /w:[ 13 1 9 0 ] /ss:0 /do:0
  and g35 (.I0(RegWr), .I1(clk), .Z(w0));   //: @(93,381) /sn:0 /delay:" 1" /w:[ 1 0 31 ]
  demux g9 (.I(SD), .E(w21), .Z0(!w8), .Z1(!w3), .Z2(!w14), .Z3(!w7), .Z4(!w15), .Z5(!w20), .Z6(!w12), .Z7(!w10));   //: @(852,169) /sn:0 /w:[ 1 0 1 0 1 1 1 0 1 1 ]
  register R4 (.Q(R4a0), .D(DIN), .EN(w15), .CLR(w4), .CK(!w0));   //: @(531,358) /w:[ 0 35 0 13 25 ]
  //: joint g7 (R10) @(532, 600) /w:[ 2 -1 1 4 ]
  or g56 (.I0(w20), .I1(Pop), .Z(w19));   //: @(746,437) /sn:0 /R:3 /w:[ 1 7 1 ]
  //: joint g58 (Pop) @(744, 301) /w:[ -1 3 4 6 ]
  //: joint g22 (w4) @(586, 337) /w:[ 5 -1 6 12 ]
  //: joint g31 (w4) @(863, 417) /w:[ 17 -1 18 28 ]
  //: joint g59 (w0) @(637, 381) /w:[ 20 22 19 -1 ]
  register R1 (.Q(R2), .D(DIN), .EN(w3), .CLR(w4), .CK(!w0));   //: @(262,449) /w:[ 7 29 1 23 11 ]
  register R3 (.Q(R3), .D(DIN), .EN(w7), .CLR(w4), .CK(!w0));   //: @(433,446) /w:[ 3 33 0 25 7 ]
  //: joint g33 (w4) @(673, 417) /w:[ 19 -1 20 26 ]
  //: joint g41 (DIN) @(717, 320) /w:[ 4 -1 3 18 ]
  //: joint g36 (w4) @(904, 337) /w:[ 1 -1 2 16 ]
  //: joint g45 (R4a0) @(531, 429) /w:[ 2 1 -1 4 ]
  //: joint g54 (DIN) @(917, 367) /w:[ 8 -1 7 14 ]
  //: joint g40 (DIN) @(433, 320) /w:[ 21 -1 22 32 ]
  //: joint g42 (DIN) @(807, 367) /w:[ 6 5 -1 16 ]
  led g52 (.I(w1));   //: @(946,591) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: joint g12 (w0) @(479, 381) /w:[ 18 24 17 -1 ]
  //: input g28 (clr) @(1034,337) /sn:0 /R:2 /w:[ 1 ]
  //: input g34 (clk) @(53,398) /sn:0 /w:[ 1 ]
  add g46 (.A(w2), .B(DIN), .S(w9), .CI(w13), .CO(w1));   //: @(949,524) /sn:0 /R:1 /w:[ 1 15 0 0 1 ]
  //: joint g57 (Pop) @(949, 297) /w:[ -1 1 2 8 ]
  mux g14 (.I0(R0t1), .I1(R2), .I2(R4), .I3(R3), .I4(R4a0), .I5(R5a1), .I6(R10), .I7(R7), .S(SA), .Z(AOUT));   //: @(279,657) /sn:0 /w:[ 9 0 5 5 7 0 0 3 0 0 ] /ss:0 /do:0
  //: input g5 (RegWr) @(46,363) /sn:0 /w:[ 0 ]
  //: joint g11 (w0) @(293, 381) /w:[ 16 26 15 -1 ]
  //: joint g21 (w4) @(388, 337) /w:[ 7 -1 8 10 ]
  //: joint g19 (R0t1) @(255, 523) /w:[ 1 -1 2 8 ]
  //: joint g61 (w0) @(542, 481) /w:[ 2 1 4 -1 ]
  //: input g20 (SD) @(780,138) /sn:0 /w:[ 0 ]
  //: joint g32 (w4) @(487, 417) /w:[ 21 -1 22 24 ]
  register R0 (.Q(R0t1), .D(DIN), .EN(w8), .CLR(w4), .CK(!w0));   //: @(181,362) /w:[ 5 27 0 9 29 ]
  led g38 (.I(R5a1));   //: @(770,677) /sn:0 /w:[ 5 ] /type:2
  //: input g0 (DIN) @(531,267) /sn:0 /R:3 /w:[ 0 ]
  //: joint g15 (R5a1) @(527, 586) /w:[ 2 -1 1 8 ]
  //: joint g43 (R2) @(262, 500) /w:[ -1 6 8 5 ]
  led t0 (.I(R0t1));   //: @(119,283) /w:[ 7 ] /type:2
  //: joint g27 (w0) @(125, 381) /w:[ 14 28 30 13 ]
  //: joint g48 (R0t1) @(181, 417) /w:[ -1 4 6 3 ]
  //: joint g62 (R5a1) @(629, 537) /w:[ 4 6 -1 3 ]
  led g37 (.I(R2));   //: @(53,495) /sn:0 /w:[ 9 ] /type:2
  and g55 (.I0(w0), .I1(Pop), .Z(w16));   //: @(648,296) /sn:0 /R:2 /w:[ 23 5 0 ]
  mux g13 (.I0(R0t1), .I1(R2), .I2(R4), .I3(R3), .I4(R4a0), .I5(R5a1), .I6(R10), .I7(R7), .S(SB), .Z(BOUT));   //: @(516,659) /sn:0 /w:[ 0 3 3 0 9 9 5 5 1 1 ] /ss:0 /do:0
  //: supply0 g53 (w13) @(947,463) /sn:0 /R:2 /w:[ 1 ]

endmodule

module ALU(Zero_signal, B, ALU_operation, A, ALU_result);
//: interface  /sz:(127, 166) /bd:[ Ti0>ALU_operation[3:0](64/127) Li0>A[31:0](46/166) Li1>B[31:0](108/166) Ro0<Zero(52/166) Ro1<ALU_result[31:0](106/166) ]
input [31:0] B;    //: /sn:0 {0}(705,303)(657,303)(657,288)(647,288){1}
//: {2}(645,286)(645,270)(598,270){3}
//: {4}(594,270)(472,270){5}
//: {6}(470,268)(470,207)(471,207){7}
//: {8}(468,270)(415,270){9}
//: {10}(596,272)(596,392)(718,392){11}
//: {12}(645,290)(645,370)(720,370){13}
supply0 w7;    //: /sn:0 {0}(669,108)(669,129)(670,129)(670,139){1}
output [31:0] ALU_result;    //: /sn:0 /dp:1 {0}(1029,324)(1108,324){1}
//: {2}(1112,324)(1147,324)(1147,292)(1194,292){3}
//: {4}(1110,326)(1110,363)(1134,363){5}
input [31:0] A;    //: /sn:0 {0}(705,279)(673,279)(673,278)(663,278){1}
//: {2}(661,276)(661,238)(614,238){3}
//: {4}(612,236)(612,149)(643,149){5}
//: {6}(610,238)(412,238){7}
//: {8}(612,240)(612,387)(718,387){9}
//: {10}(661,280)(661,365)(720,365){11}
supply0 w0;    //: /sn:0 {0}(729,225)(729,250)(730,250)(730,260){1}
supply0 w3;    //: /sn:0 {0}(554,108)(554,134)(555,134)(555,144){1}
supply0 [31:0] w20;    //: /sn:0 {0}(805,115)(805,119)(899,119){1}
input [3:0] ALU_operation;    //: /sn:0 {0}(428,544)(723,544)(723,543)(1016,543){1}
//: {2}(1017,543)(1078,543){3}
output Zero_signal;    //: /sn:0 /dp:1 {0}(1219,391)(1342,391)(1342,388)(1352,388){1}
supply0 [31:0] w5;    //: /sn:0 {0}(825,318)(857,318)(857,317)(867,317){1}
//: {2}(869,315)(869,314)(1000,314){3}
//: {4}(869,319)(869,320)(983,320){5}
//: {6}(987,320)(1000,320){7}
//: {8}(985,322)(985,327)(1000,327){9}
wire [31:0] w16;    //: /sn:0 /dp:3 {0}(1000,307)(818,307)(818,160){1}
//: {2}(818,159)(818,149)(803,149)(803,161)(686,161){3}
wire [31:0] w13;    //: /sn:0 {0}(527,156)(515,156)(515,155){1}
//: {2}(517,153)(522,153)(522,99)(899,99){3}
//: {4}(513,153)(465,153)(465,133){5}
wire Zero;    //: /sn:0 /dp:1 {0}(822,160)(915,160)(915,132){1}
wire [31:0] w22;    //: /sn:0 /dp:1 {0}(582,170)(628,170)(628,168)(643,168){1}
wire [31:0] w18;    //: /sn:0 {0}(741,368)(793,368)(793,347)(1000,347){1}
wire [31:0] w12;    //: /sn:0 {0}(487,207)(500,207)(500,178)(527,178){1}
wire w19;    //: /sn:0 /dp:1 {0}(688,218)(688,193)(666,193)(666,183){1}
wire [2:0] w10;    //: /sn:0 {0}(1017,538)(1017,442)(1016,442)(1016,347){1}
wire w21;    //: /sn:0 {0}(556,196)(556,215)(569,215)(569,225){1}
wire [31:0] w17;    //: /sn:0 {0}(928,109)(990,109)(990,300)(1000,300){1}
wire w14;    //: /sn:0 {0}(1155,363)(1193,363)(1193,391)(1203,391){1}
wire w11;    //: /sn:0 {0}(731,316)(731,326)(754,326)(754,345){1}
wire [31:0] w15;    //: /sn:0 {0}(753,288)(800,288)(800,334)(1000,334){1}
wire [31:0] w9;    //: /sn:0 {0}(739,390)(803,390)(803,340)(1000,340){1}
//: enddecls

  or g4 (.I0(A), .I1(B), .Z(w9));   //: @(729,390) /sn:0 /w:[ 9 11 0 ]
  //: joint g8 (A) @(612, 238) /w:[ 3 4 6 8 ]
  and g3 (.I0(A), .I1(B), .Z(w18));   //: @(731,368) /sn:0 /w:[ 11 13 0 ]
  //: supply0 g16 (w5) @(819,318) /sn:0 /R:3 /w:[ 0 ]
  not g17 (.I(w14), .Z(Zero_signal));   //: @(1209,391) /sn:0 /w:[ 1 0 ]
  CLA32 g26 (.Cin(w7), .A(A), .B(w22), .Cout(w19), .S(w16));   //: @(644, 140) /sz:(41, 42) /sn:0 /p:[ Ti0>1 Li0>5 Li1>1 Bo0<1 Ro0<3 ]
  or g2 (.I0(ALU_result), .Z(w14));   //: @(1145,363) /sn:0 /w:[ 5 0 ]
  //: joint g23 (B) @(470, 270) /w:[ 5 6 8 -1 ]
  //: joint g30 (w5) @(869, 317) /w:[ -1 2 1 4 ]
  //: supply0 g24 (w3) @(554,102) /sn:0 /R:2 /w:[ 0 ]
  //: joint g1 (B) @(645, 288) /w:[ 1 2 -1 12 ]
  mux g29 (.I0(w18), .I1(w9), .I2(w15), .I3(w5), .I4(w5), .I5(w5), .I6(w16), .I7(w17), .S(w10), .Z(ALU_result));   //: @(1016,324) /sn:0 /R:1 /w:[ 1 1 1 9 7 3 0 1 1 0 ] /ss:0 /do:0
  //: output g18 (Zero_signal) @(1349,388) /sn:0 /w:[ 1 ]
  //: supply0 g10 (w0) @(729,219) /sn:0 /R:2 /w:[ 0 ]
  led g25 (.I(w21));   //: @(569,232) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: input g6 (B) @(413,270) /sn:0 /w:[ 9 ]
  //: joint g9 (B) @(596, 270) /w:[ 3 -1 4 10 ]
  //: joint g7 (A) @(661, 278) /w:[ 1 2 -1 10 ]
  //: joint g31 (w5) @(985, 320) /w:[ 6 -1 5 8 ]
  //: joint g22 (w13) @(515, 153) /w:[ 2 -1 4 1 ]
  tran g33(.Z(Zero), .I(w16[31]));   //: @(816,160) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  //: input g12 (ALU_operation) @(426,544) /sn:0 /w:[ 0 ]
  led g28 (.I(w19));   //: @(688,225) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: supply0 g34 (w20) @(805,109) /sn:0 /R:2 /w:[ 0 ]
  //: input g5 (A) @(410,238) /sn:0 /w:[ 7 ]
  led g11 (.I(w11));   //: @(754,352) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: output g14 (ALU_result) @(1191,292) /sn:0 /w:[ 3 ]
  //: dip g21 (w13) @(465,123) /sn:0 /w:[ 5 ] /st:1
  CLA32 g19 (.Cin(w3), .A(w13), .B(w12), .Cout(w21), .S(w22));   //: @(528, 145) /sz:(53, 50) /sn:0 /p:[ Ti0>1 Li0>0 Li1>1 Bo0<0 Ro0<0 ]
  not g20 (.I(B), .Z(w12));   //: @(477,207) /sn:0 /w:[ 7 0 ]
  mux g32 (.I0(w20), .I1(w13), .S(Zero), .Z(w17));   //: @(915,109) /sn:0 /R:1 /w:[ 1 3 1 0 ] /ss:0 /do:0
  //: joint g15 (ALU_result) @(1110, 324) /w:[ 2 -1 1 4 ]
  CLA32 g0 (.Cin(w0), .A(B), .B(A), .Cout(w11), .S(w15));   //: @(706, 261) /sz:(46, 54) /sn:0 /p:[ Ti0>1 Li0>0 Li1>0 Bo0<0 Ro0<0 ]
  //: supply0 g27 (w7) @(669,102) /sn:0 /R:2 /w:[ 0 ]
  tran g13(.Z(w10), .I(ALU_operation[2:0]));   //: @(1017,541) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0

endmodule

module EXE(ALU_result, Zero_signal, data_read_2, data_read_1, INM32, PCNext, branch_target, ALU_operation);
//: interface  /sz:(185, 314) /bd:[ Ti0>ALU_operation[3:0](85/185) Li0>data_read_2[31:0](272/314) Li1>data_read_1[31:0](239/314) Li2>PCNext[31:0](91/314) Li3>INM32[31:0](126/314) Ro0<Zero_signal(242/314) Ro1<ALU_result[31:0](283/314) Ro2<branch_target[31:0](90/314) ]
output [31:0] ALU_result;    //: /sn:0 {0}(540,374)(679,374){1}
input [3:0] ALU_operation;    //: /sn:0 {0}(406,120)(464,120)(464,244){1}
input [31:0] data_read_2;    //: /sn:0 {0}(166,377)(387,377){1}
input [31:0] PCNext;    //: /sn:0 {0}(113,514)(447,514)(447,559)(455,559){1}
output Zero_signal;    //: /sn:0 {0}(540,308)(675,308){1}
output [31:0] branch_target;    //: /sn:0 /dp:1 {0}(543,582)(593,582)(593,572)(615,572){1}
input [31:0] INM32;    //: /sn:0 /dp:1 {0}(116,623)(447,623)(447,596)(455,596){1}
supply0 w5;    //: /sn:0 {0}(499,510)(499,529)(501,529)(501,539){1}
input [31:0] data_read_1;    //: /sn:0 {0}(170,301)(387,301){1}
wire w4;    //: /sn:0 {0}(502,625)(502,670){1}
//: enddecls

  led g8 (.I(w4));   //: @(502,677) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: output g4 (ALU_result) @(676,374) /sn:0 /w:[ 1 ]
  //: output g3 (Zero_signal) @(672,308) /sn:0 /w:[ 1 ]
  //: input g2 (data_read_2) @(164,377) /sn:0 /w:[ 0 ]
  //: input g1 (data_read_1) @(168,301) /sn:0 /w:[ 0 ]
  //: input g10 (INM32) @(114,623) /sn:0 /w:[ 0 ]
  //: input g9 (PCNext) @(111,514) /sn:0 /w:[ 0 ]
  //: supply0 g7 (w5) @(499,504) /sn:0 /R:2 /w:[ 0 ]
  CLA32 g12 (.Cin(w5), .A(PCNext), .B(INM32), .Cout(w4), .S(branch_target));   //: @(456, 540) /sz:(86, 84) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Bo0<0 Ro0<0 ]
  //: output g11 (branch_target) @(612,572) /sn:0 /w:[ 1 ]
  //: input g5 (ALU_operation) @(404,120) /sn:0 /w:[ 0 ]
  ALU g0 (.ALU_operation(ALU_operation), .B(data_read_2), .A(data_read_1), .ALU_result(ALU_result), .Zero_signal(Zero_signal));   //: @(388, 245) /sz:(151, 203) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Ro0<0 Ro1<0 ]

endmodule

module BRegs32x32(Read2, Write, Read1, Data2, Data1, clr, Pop, clk, RegWrite, WriteData);
//: interface  /sz:(147, 182) /bd:[ Ti0>clr(66/147) Ti1>clr(66/147) Ti2>Pop(105/147) Ti3>clr(66/147) Li0>WriteData[31:0](148/182) Li1>Write[4:0](108/182) Li2>Read2[4:0](72/182) Li3>Read1[4:0](32/182) Li4>WriteData[31:0](148/182) Li5>Write[4:0](108/182) Li6>Read2[4:0](72/182) Li7>Read1[4:0](32/182) Li8>Read1[4:0](32/182) Li9>Read2[4:0](72/182) Li10>Write[4:0](108/182) Li11>WriteData[31:0](148/182) Bi0>RegWrite(40/147) Bi1>clk(108/147) Bi2>RegWrite(40/147) Bi3>clk(108/147) Bi4>clk(108/147) Bi5>RegWrite(40/147) Ro0<Data2[31:0](139/182) Ro1<Data1[31:0](47/182) Ro2<Data2[31:0](139/182) Ro3<Data1[31:0](47/182) Ro4<Data1[31:0](47/182) Ro5<Data2[31:0](139/182) ]
output [31:0] Data2;    //: /sn:0 {0}(668,485)(668,472)(669,472)(669,445){1}
input Pop;    //: /sn:0 {0}(863,67)(708,67)(708,157){1}
input [4:0] Write;    //: /sn:0 {0}(-238,-38)(-138,-38)(-138,-37)(-66,-37){1}
//: {2}(-65,-37)(-28,-37){3}
//: {4}(-27,-37)(-16,-37){5}
input [31:0] WriteData;    //: /sn:0 {0}(670,157)(670,75)(481,75){1}
//: {2}(477,75)(292,75){3}
//: {4}(288,75)(89,75){5}
//: {6}(85,75)(-104,75)(-104,73)(-237,73){7}
//: {8}(87,77)(87,157){9}
//: {10}(290,77)(290,107)(291,107)(291,152){11}
//: {12}(479,77)(479,117)(478,117)(478,157){13}
supply1 w21;    //: /sn:0 {0}(82,3)(57,3)(57,-11){1}
output [31:0] Data1;    //: /sn:0 {0}(59,382)(59,465){1}
input RegWrite;    //: /sn:0 {0}(-237,263)(-71,263){1}
//: {2}(-67,263)(171,263){3}
//: {4}(175,263)(370,263){5}
//: {6}(374,263)(552,263)(552,219)(556,219){7}
//: {8}(372,261)(372,219)(383,219){9}
//: {10}(173,261)(173,214)(183,214){11}
//: {12}(-69,261)(-69,219)(-38,219){13}
input clr;    //: /sn:0 {0}(722,193)(732,193)(732,-83)(543,-83){1}
//: {2}(539,-83)(355,-83){3}
//: {4}(351,-83)(150,-83){5}
//: {6}(146,-83)(-44,-83)(-44,-92)(-235,-92){7}
//: {8}(148,-81)(148,193)(139,193){9}
//: {10}(353,-81)(353,188)(343,188){11}
//: {12}(541,-81)(541,193)(530,193){13}
input clk;    //: /sn:0 {0}(556,214)(542,214)(542,285)(364,285){1}
//: {2}(362,283)(362,214)(383,214){3}
//: {4}(360,285)(167,285){5}
//: {6}(165,283)(165,209)(183,209){7}
//: {8}(163,285)(-56,285){9}
//: {10}(-58,283)(-58,214)(-38,214){11}
//: {12}(-60,285)(-237,285){13}
input [4:0] Read1;    //: {0}(-237,96)(-208,96)(-208,95)(-124,95){1}
//: {2}(-123,95)(-96,95){3}
//: {4}(-95,95)(-78,95){5}
input [4:0] Read2;    //: {0}(-237,145)(-141,145){1}
//: {2}(-140,145)(-123,145)(-123,144)(-94,144){3}
//: {4}(-93,144)(-79,144){5}
wire w16;    //: /sn:0 {0}(39,205)(-50,205)(-50,39)(88,39)(88,19){1}
wire [1:0] w6;    //: /sn:0 {0}(36,369)(-123,369)(-123,99){1}
wire w4;    //: /sn:0 {0}(112,19)(112,46)(369,46)(369,205)(430,205){1}
wire w22;    //: /sn:0 {0}(404,217)(430,217){1}
wire [31:0] w0;    //: /sn:0 {0}(651,416)(651,398)(105,398)(105,228){1}
wire [31:0] R2;    //: {0}(65,353)(65,319)(468,319)(468,228){1}
wire [31:0] w3;    //: /sn:0 {0}(77,353)(77,334)(660,334)(660,228){1}
wire w20;    //: /sn:0 {0}(124,19)(124,29)(557,29)(557,205)(622,205){1}
wire [2:0] w18;    //: /sn:0 {0}(430,180)(402,180)(402,125){1}
//: {2}(404,123)(590,123)(590,180)(622,180){3}
//: {4}(400,123)(279,123)(279,122)(212,122){5}
//: {6}(208,122)(8,122){7}
//: {8}(4,122)(-93,122)(-93,139){9}
//: {10}(6,124)(6,180)(39,180){11}
//: {12}(210,124)(210,175)(243,175){13}
wire [2:0] w19;    //: /sn:0 {0}(430,169)(419,169)(419,109){1}
//: {2}(421,107)(607,107)(607,169)(622,169){3}
//: {4}(417,107)(297,107)(297,106)(231,106){5}
//: {6}(227,106)(25,106){7}
//: {8}(21,106)(-95,106)(-95,99){9}
//: {10}(23,108)(23,169)(39,169){11}
//: {12}(229,108)(229,164)(243,164){13}
wire [1:0] w10;    //: /sn:0 {0}(-140,149)(-140,432)(646,432){1}
wire w23;    //: /sn:0 {0}(577,217)(622,217){1}
wire [2:0] w24;    //: /sn:0 {0}(430,193)(381,193)(381,141){1}
//: {2}(383,139)(569,139)(569,193)(622,193){3}
//: {4}(379,139)(260,139)(260,138)(195,138){5}
//: {6}(191,138)(-13,138){7}
//: {8}(-17,138)(-65,138)(-65,-33){9}
//: {10}(-15,140)(-15,193)(39,193){11}
//: {12}(193,140)(193,188)(243,188){13}
wire w1;    //: /sn:0 {0}(-17,217)(39,217){1}
wire w31;    //: /sn:0 {0}(243,200)(178,200)(178,60)(100,60)(100,19){1}
wire [31:0] R3;    //: {0}(688,228)(688,322)(687,322)(687,416){1}
wire [31:0] R1;    //: {0}(281,223)(281,308)(53,308)(53,353){1}
wire w2;    //: /sn:0 {0}(243,212)(204,212){1}
wire [1:0] w11;    //: /sn:0 {0}(-27,-33)(-27,-23)(106,-23)(106,-10){1}
wire [31:0] R0;    //: {0}(77,228)(77,299)(41,299)(41,353){1}
wire [31:0] w5;    //: /sn:0 {0}(675,416)(675,372)(496,372)(496,228){1}
wire [31:0] w9;    //: /sn:0 {0}(663,416)(663,387)(309,387)(309,223){1}
//: enddecls

  //: joint g44 (clr) @(353, -83) /w:[ 3 -1 4 10 ]
  //: input g4 (Read2) @(-239,145) /sn:0 /w:[ 0 ]
  //: joint g8 (w18) @(6, 122) /w:[ 7 -1 8 10 ]
  //: joint g47 (clr) @(541, -83) /w:[ 1 -1 2 12 ]
  //: joint g16 (clk) @(165, 285) /w:[ 5 6 8 -1 ]
  //: input g3 (Write) @(-240,-38) /sn:0 /w:[ 0 ]
  //: joint g26 (w19) @(229, 106) /w:[ 5 -1 6 12 ]
  //: input g17 (Read1) @(-239,96) /sn:0 /w:[ 0 ]
  //: output g2 (Data2) @(668,482) /sn:0 /R:3 /w:[ 0 ]
  tran g30(.Z(w10), .I(Read2[4:3]));   //: @(-140,143) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g23(.Z(w24), .I(Write[2:0]));   //: @(-65,-39) /sn:0 /R:1 /w:[ 9 1 2 ] /ss:1
  Regs8x32 g24 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w31), .clk(w2), .clr(clr), .AOUT(R1), .BOUT(w9));   //: @(244, 153) /sz:(98, 69) /sn:0 /p:[ Ti0>11 Li0>13 Li1>13 Li2>13 Li3>0 Li4>0 Ri0>11 Bo0<0 Bo1<1 ]
  //: joint g39 (RegWrite) @(372, 263) /w:[ 6 8 5 -1 ]
  //: output g1 (Data1) @(59,462) /sn:0 /R:3 /w:[ 1 ]
  Regs8x32 g29 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w4), .clk(w22), .clr(clr), .AOUT(R2), .BOUT(w5));   //: @(431, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>13 Li0>0 Li1>0 Li2>0 Li3>1 Li4>1 Ri0>13 Bo0<1 Bo1<1 ]
  //: comment g51 /dolink:0 /link:"" @(395,229) /sn:0
  //: /line:"Regs 16-23"
  //: /end
  tran g18(.Z(w19), .I(Read1[2:0]));   //: @(-95,93) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:1
  //: joint g25 (w18) @(210, 122) /w:[ 5 -1 6 12 ]
  //: supply1 g10 (w21) @(68,-11) /sn:0 /w:[ 1 ]
  //: comment g49 /dolink:0 /link:"" @(210,225) /sn:0
  //: /line:"Regs 8-15"
  //: /end
  Regs8x32 g6 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w16), .clk(w1), .clr(clr), .AOUT(R0), .BOUT(w0));   //: @(40, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>9 Li0>11 Li1>11 Li2>11 Li3>0 Li4>1 Ri0>9 Bo0<0 Bo1<1 ]
  //: comment g50 /dolink:0 /link:"" @(585,229) /sn:0
  //: /line:"Regs 24-31"
  //: /end
  and g35 (.I0(clk), .I1(RegWrite), .Z(w22));   //: @(394,217) /sn:0 /delay:" 1" /w:[ 3 9 0 ]
  demux g9 (.I(w11), .E(w21), .Z0(w16), .Z1(w31), .Z2(w4), .Z3(w20));   //: @(106,3) /sn:0 /w:[ 1 0 1 1 0 0 ]
  //: joint g7 (w19) @(23, 106) /w:[ 7 -1 8 10 ]
  tran g22(.Z(w18), .I(Read2[2:0]));   //: @(-93,142) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:0
  tran g31(.Z(w6), .I(Read1[4:3]));   //: @(-123,93) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  and g33 (.I0(clk), .I1(RegWrite), .Z(w1));   //: @(-27,217) /sn:0 /delay:" 1" /w:[ 11 13 0 ]
  //: joint g45 (WriteData) @(479, 75) /w:[ 1 -1 2 12 ]
  //: joint g41 (w19) @(419, 107) /w:[ 2 -1 4 1 ]
  and g36 (.I0(clk), .I1(RegWrite), .Z(w23));   //: @(567,217) /sn:0 /delay:" 1" /w:[ 0 7 0 ]
  //: joint g40 (w18) @(402, 123) /w:[ 2 -1 4 1 ]
  //: input g42 (clr) @(-237,-92) /sn:0 /w:[ 7 ]
  //: input g52 (Pop) @(865,67) /sn:0 /R:2 /w:[ 0 ]
  //: input g12 (clk) @(-239,285) /sn:0 /w:[ 13 ]
  Regs8x324 g46 (.Pop(Pop), .DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w20), .clk(w23), .clr(clr), .AOUT(w3), .BOUT(R3));   //: @(623, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>3 Li1>3 Li2>3 Li3>1 Li4>1 Ri0>0 Bo0<1 Bo1<0 ]
  //: joint g28 (w24) @(381, 139) /w:[ 2 -1 4 1 ]
  and g34 (.I0(clk), .I1(RegWrite), .Z(w2));   //: @(194,212) /sn:0 /delay:" 1" /w:[ 7 11 1 ]
  tran g5(.Z(w11), .I(Write[4:3]));   //: @(-27,-39) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  mux g14 (.I0(R0), .I1(R1), .I2(R2), .I3(w3), .S(w6), .Z(Data1));   //: @(59,369) /sn:0 /w:[ 1 1 0 0 0 0 ] /ss:0 /do:0
  //: joint g11 (w24) @(-15, 138) /w:[ 7 -1 8 10 ]
  //: joint g21 (w24) @(193, 138) /w:[ 5 -1 6 12 ]
  //: joint g19 (clk) @(-58, 285) /w:[ 9 10 12 -1 ]
  //: joint g20 (WriteData) @(87, 75) /w:[ 5 -1 6 8 ]
  //: input g32 (RegWrite) @(-239,263) /sn:0 /w:[ 0 ]
  //: input g0 (WriteData) @(-239,73) /sn:0 /w:[ 7 ]
  //: joint g43 (clr) @(148, -83) /w:[ 5 -1 6 8 ]
  //: joint g15 (clk) @(362, 285) /w:[ 1 2 4 -1 ]
  //: joint g38 (RegWrite) @(173, 263) /w:[ 4 10 3 -1 ]
  //: comment g48 /dolink:0 /link:"" @(11,228) /sn:0
  //: /line:"Regs 0-7"
  //: /end
  //: joint g27 (WriteData) @(290, 75) /w:[ 3 -1 4 10 ]
  //: joint g37 (RegWrite) @(-69, 263) /w:[ 2 12 1 -1 ]
  mux g13 (.I0(w0), .I1(w9), .I2(w5), .I3(R3), .S(w10), .Z(Data2));   //: @(669,432) /sn:0 /w:[ 0 0 0 1 1 1 ] /ss:0 /do:0

endmodule

module Regs8x32(SB, SA, BOUT, AOUT, clr, clk, RegWr, SD, DIN);
//: interface  /sz:(98, 69) /bd:[ Ti0>DIN[31:0](47/98) Li0>SD[2:0](35/69) Li1>SA[2:0](11/69) Li2>SB[2:0](22/69) Li3>RegWr(47/69) Li4>clk(59/69) Ri0>clr(35/69) Bo0<AOUT[31:0](37/98) Bo1<BOUT[31:0](65/98) ]
input [31:0] DIN;    //: /sn:0 {0}(181,352)(181,320)(260,320){1}
//: {2}(264,320)(338,320){3}
//: {4}(342,320)(431,320){5}
//: {6}(435,320)(529,320){7}
//: {8}(533,320)(627,320){9}
//: {10}(631,320)(715,320){11}
//: {12}(719,320)(807,320)(807,429){13}
//: {14}(717,322)(717,352){15}
//: {16}(629,322)(629,433){17}
//: {18}(531,318)(531,269){19}
//: {20}(531,322)(531,348){21}
//: {22}(433,322)(433,436){23}
//: {24}(340,322)(340,351){25}
//: {26}(262,322)(262,439){27}
output [31:0] BOUT;    //: /sn:0 {0}(516,697)(516,672){1}
input [2:0] SD;    //: /sn:0 {0}(782,138)(852,138)(852,156){1}
input [2:0] SB;    //: /sn:0 {0}(466,659)(493,659){1}
supply1 w21;    //: /sn:0 {0}(828,169)(801,169)(801,153){1}
input RegWr;    //: /sn:0 {0}(48,363)(68,363)(68,378)(82,378){1}
input clr;    //: /sn:0 /dp:1 {0}(959,337)(1032,337){1}
input [2:0] SA;    //: /sn:0 {0}(256,657)(231,657){1}
input clk;    //: /sn:0 {0}(82,383)(68,383)(68,398)(55,398){1}
output [31:0] AOUT;    //: /sn:0 {0}(279,670)(279,702){1}
wire [31:0] w16;    //: /sn:0 {0}(531,369)(531,435){1}
//: {2}(533,437)(581,437)(581,177){3}
//: {4}(531,439)(531,574)(520,574){5}
//: {6}(516,574)(282,574)(282,641){7}
//: {8}(518,576)(518,587)(519,587)(519,643){9}
wire w7;    //: /sn:0 {0}(472,451)(513,451)(513,405)(848,405)(848,185){1}
wire [31:0] R5;    //: {0}(288,641)(288,586)(525,586){1}
//: {2}(529,586)(629,586)(629,529){3}
//: {4}(631,527)(684,527)(684,290){5}
//: {6}(629,525)(629,454){7}
//: {8}(527,588)(527,617)(525,617)(525,643){9}
wire w4;    //: /sn:0 {0}(943,337)(906,337){1}
//: {2}(902,337)(767,337){3}
//: {4}(763,337)(588,337){5}
//: {6}(584,337)(390,337){7}
//: {8}(386,337)(231,337)(231,357)(220,357){9}
//: {10}(388,339)(388,356)(379,356){11}
//: {12}(586,339)(586,353)(570,353){13}
//: {14}(765,339)(765,357)(756,357){15}
//: {16}(904,339)(904,417)(865,417){17}
//: {18}(861,417)(675,417){19}
//: {20}(671,417)(489,417){21}
//: {22}(485,417)(302,417)(302,444)(301,444){23}
//: {24}(487,419)(487,441)(472,441){25}
//: {26}(673,419)(673,438)(668,438){27}
//: {28}(863,419)(863,434)(846,434){29}
wire w3;    //: /sn:0 {0}(835,185)(835,397)(330,397)(330,454)(301,454){1}
wire w0;    //: /sn:0 {0}(770,439)(764,439)(764,481)(579,481){1}
//: {2}(577,479)(577,443)(592,443){3}
//: {4}(575,481)(390,481){5}
//: {6}(388,479)(388,446)(396,446){7}
//: {8}(386,481)(214,481){9}
//: {10}(212,479)(212,449)(225,449){11}
//: {12}(210,481)(125,481)(125,383){13}
//: {14}(127,381)(291,381){15}
//: {16}(295,381)(477,381){17}
//: {18}(481,381)(660,381)(660,362)(680,362){19}
//: {20}(479,379)(479,358)(494,358){21}
//: {22}(293,379)(293,361)(303,361){23}
//: {24}(125,379)(125,362)(144,362){25}
//: {26}(123,381)(103,381){27}
wire [31:0] R2;    //: {0}(262,641)(262,537){1}
//: {2}(264,535)(499,535)(499,643){3}
//: {4}(262,533)(262,495){5}
//: {6}(262,491)(262,460){7}
//: {8}(260,493)(44,493)(44,534){9}
wire [31:0] R7;    //: {0}(807,450)(807,569){1}
//: {2}(809,571)(951,571)(951,541){3}
//: {4}(807,573)(807,609)(541,609){5}
//: {6}(537,609)(302,609)(302,641){7}
//: {8}(539,611)(539,643){9}
wire w12;    //: /sn:0 {0}(756,367)(787,367)(787,258)(868,258)(868,185){1}
wire w10;    //: /sn:0 {0}(846,444)(875,444)(875,185){1}
wire [31:0] R4;    //: {0}(340,372)(340,408){1}
//: {2}(342,410)(373,410)(373,271){3}
//: {4}(340,412)(340,545){5}
//: {6}(342,547)(505,547)(505,643){7}
//: {8}(338,547)(268,547)(268,641){9}
wire [31:0] R3;    //: {0}(512,643)(512,559)(435,559){1}
//: {2}(433,557)(433,510){3}
//: {4}(433,506)(433,457){5}
//: {6}(431,508)(393,508)(393,707){7}
//: {8}(431,559)(275,559)(275,641){9}
wire w8;    //: /sn:0 {0}(220,367)(249,367)(249,213)(828,213)(828,185){1}
wire Z5;    //: /sn:0 {0}(861,185)(861,413)(700,413)(700,448)(668,448){1}
wire w14;    //: /sn:0 {0}(379,366)(414,366)(414,229)(841,229)(841,185){1}
wire [31:0] R0;    //: {0}(492,643)(492,523)(257,523){1}
//: {2}(253,523)(181,523)(181,423){3}
//: {4}(181,419)(181,373){5}
//: {6}(179,421)(119,421)(119,280){7}
//: {8}(255,525)(255,641){9}
wire w15;    //: /sn:0 {0}(570,363)(608,363)(608,244)(855,244)(855,185){1}
wire [31:0] R10;    //: /sn:0 {0}(295,641)(295,600)(530,600){1}
//: {2}(534,600)(717,600)(717,571){3}
//: {4}(719,569)(750,569)(750,641){5}
//: {6}(717,567)(717,373){7}
//: {8}(532,602)(532,643){9}
//: enddecls

  led g44 (.I(R5));   //: @(684,283) /sn:0 /w:[ 5 ] /type:2
  //: input g4 (SB) @(464,659) /sn:0 /w:[ 0 ]
  //: joint g8 (w16) @(518, 574) /w:[ 5 -1 6 8 ]
  led g47 (.I(R7));   //: @(951,534) /sn:0 /w:[ 3 ] /type:2
  //: joint g16 (R3) @(433, 559) /w:[ 1 2 8 -1 ]
  //: input g3 (SA) @(229,657) /sn:0 /w:[ 1 ]
  //: joint g26 (DIN) @(340, 320) /w:[ 4 -1 3 24 ]
  //: joint g17 (R4) @(340, 547) /w:[ 6 5 8 -1 ]
  //: output g2 (BOUT) @(516,694) /sn:0 /R:3 /w:[ 0 ]
  register R5 (.Q(R5), .D(DIN), .EN(Z5), .CLR(w4), .CK(!w0));   //: @(629,443) /w:[ 7 17 1 27 3 ]
  //: joint g30 (w0) @(212, 481) /w:[ 9 10 12 -1 ]
  //: joint g23 (w4) @(765, 337) /w:[ 3 -1 4 14 ]
  //: joint g24 (DIN) @(531, 320) /w:[ 8 18 7 20 ]
  //: joint g39 (DIN) @(262, 320) /w:[ 2 -1 1 26 ]
  //: output g1 (AOUT) @(279,699) /sn:0 /R:3 /w:[ 1 ]
  //: joint g29 (w0) @(388, 481) /w:[ 5 6 8 -1 ]
  //: joint g51 (R5) @(629, 527) /w:[ 4 6 -1 3 ]
  register R2 (.Q(R4), .D(DIN), .EN(w14), .CLR(w4), .CK(!w0));   //: @(340,361) /w:[ 0 25 0 11 23 ]
  //: joint g18 (R2) @(262, 535) /w:[ 2 4 -1 1 ]
  register R7 (.Q(R7), .D(DIN), .EN(w10), .CLR(w4), .CK(!w0));   //: @(807,439) /w:[ 0 13 0 29 0 ]
  not g25 (.I(clr), .Z(w4));   //: @(953,337) /sn:0 /R:2 /w:[ 0 0 ]
  //: supply1 g10 (w21) @(812,153) /sn:0 /w:[ 1 ]
  //: joint g49 (R7) @(807, 571) /w:[ 2 1 -1 4 ]
  //: joint g50 (R10) @(717, 569) /w:[ 4 6 -1 3 ]
  register R6 (.Q(R10), .D(DIN), .EN(w12), .CLR(w4), .CK(!w0));   //: @(717,362) /w:[ 7 15 0 15 19 ]
  //: joint g6 (R7) @(539, 609) /w:[ 5 -1 6 8 ]
  led g56 (.I(R3));   //: @(393,714) /sn:0 /R:2 /w:[ 7 ] /type:2
  and g35 (.I0(RegWr), .I1(clk), .Z(w0));   //: @(93,381) /sn:0 /delay:" 1" /w:[ 1 0 27 ]
  demux g9 (.I(SD), .E(w21), .Z0(!w8), .Z1(!w3), .Z2(!w14), .Z3(!w7), .Z4(!w15), .Z5(!Z5), .Z6(!w12), .Z7(!w10));   //: @(852,169) /sn:0 /w:[ 1 0 1 0 1 1 1 0 1 1 ]
  register R4 (.Q(w16), .D(DIN), .EN(w15), .CLR(w4), .CK(!w0));   //: @(531,358) /w:[ 0 21 0 13 21 ]
  //: joint g7 (R10) @(532, 600) /w:[ 2 -1 1 8 ]
  //: joint g22 (w4) @(586, 337) /w:[ 5 -1 6 12 ]
  //: joint g31 (w4) @(863, 417) /w:[ 17 -1 18 28 ]
  register R1 (.Q(R2), .D(DIN), .EN(w3), .CLR(w4), .CK(!w0));   //: @(262,449) /w:[ 7 27 1 23 11 ]
  register R3 (.Q(R3), .D(DIN), .EN(w7), .CLR(w4), .CK(!w0));   //: @(433,446) /w:[ 5 23 0 25 7 ]
  led g54 (.I(R2));   //: @(44,541) /sn:0 /R:2 /w:[ 9 ] /type:2
  led g45 (.I(R10));   //: @(750,648) /sn:0 /R:2 /w:[ 5 ] /type:2
  //: joint g33 (w4) @(673, 417) /w:[ 19 -1 20 26 ]
  //: joint g41 (DIN) @(717, 320) /w:[ 12 -1 11 14 ]
  //: joint g36 (w4) @(904, 337) /w:[ 1 -1 2 16 ]
  //: joint g52 (R4) @(340, 410) /w:[ 2 1 -1 4 ]
  //: joint g40 (DIN) @(433, 320) /w:[ 6 -1 5 22 ]
  //: joint g42 (DIN) @(629, 320) /w:[ 10 -1 9 16 ]
  //: joint g12 (w0) @(479, 381) /w:[ 18 20 17 -1 ]
  //: joint g57 (R3) @(433, 508) /w:[ -1 4 6 3 ]
  led g46 (.I(w16));   //: @(581,170) /sn:0 /w:[ 3 ] /type:2
  //: input g28 (clr) @(1034,337) /sn:0 /R:2 /w:[ 1 ]
  //: input g34 (clk) @(53,398) /sn:0 /w:[ 1 ]
  mux g14 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SA), .Z(AOUT));   //: @(279,657) /sn:0 /w:[ 9 0 9 9 7 0 0 7 0 0 ] /ss:0 /do:0
  //: input g5 (RegWr) @(46,363) /sn:0 /w:[ 0 ]
  //: joint g11 (w0) @(293, 381) /w:[ 16 22 15 -1 ]
  //: joint g21 (w4) @(388, 337) /w:[ 7 -1 8 10 ]
  //: joint g19 (R0) @(255, 523) /w:[ 1 -1 2 8 ]
  //: input g20 (SD) @(780,138) /sn:0 /w:[ 0 ]
  //: joint g32 (w4) @(487, 417) /w:[ 21 -1 22 24 ]
  register R0 (.Q(R0), .D(DIN), .EN(w8), .CLR(w4), .CK(!w0));   //: @(181,362) /w:[ 5 0 0 9 25 ]
  led g43 (.I(R4));   //: @(373,264) /sn:0 /w:[ 3 ] /type:2
  //: input g0 (DIN) @(531,267) /sn:0 /R:3 /w:[ 19 ]
  //: joint g15 (R5) @(527, 586) /w:[ 2 -1 1 8 ]
  //: joint g38 (w0) @(577, 481) /w:[ 1 2 4 -1 ]
  //: joint g48 (R0) @(181, 421) /w:[ -1 4 6 3 ]
  //: joint g27 (w0) @(125, 381) /w:[ 14 24 26 13 ]
  led g37 (.I(R0));   //: @(119,273) /sn:0 /w:[ 7 ] /type:2
  //: joint g55 (R2) @(262, 493) /w:[ -1 6 8 5 ]
  //: joint g53 (w16) @(531, 437) /w:[ 2 1 -1 4 ]
  mux g13 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SB), .Z(BOUT));   //: @(516,659) /sn:0 /w:[ 0 3 7 0 9 9 9 9 1 1 ] /ss:0 /do:0

endmodule

module FA(Cout, S, Cin, B, A);
//: interface  /sz:(40, 40) /bd:[ Ti0>Cin(19/40) Li0>B(29/40) Li1>A(13/40) Ro0<Cout(32/40) Ro1<S(15/40) ]
input B;    //: /sn:0 {0}(160,154)(128,154)(128,104)(115,104){1}
//: {2}(113,102)(113,91)(123,91){3}
//: {4}(111,104)(95,104){5}
input A;    //: /sn:0 {0}(97,85)(102,85){1}
//: {2}(106,85)(113,85)(113,86)(123,86){3}
//: {4}(104,87)(104,159)(160,159){5}
input Cin;    //: /sn:0 {0}(99,123)(154,123){1}
//: {2}(156,121)(156,100)(170,100){3}
//: {4}(156,125)(156,129)(160,129){5}
output Cout;    //: /sn:0 {0}(277,142)(233,142){1}
output S;    //: /sn:0 {0}(275,100)(201,100)(201,98)(191,98){1}
wire w13;    //: /sn:0 /dp:1 {0}(212,144)(191,144)(191,157)(181,157){1}
wire w7;    //: /sn:0 {0}(160,134)(149,134)(149,91){1}
//: {2}(151,89)(153,89)(153,95)(170,95){3}
//: {4}(147,89)(144,89){5}
wire w12;    //: /sn:0 /dp:1 {0}(212,139)(191,139)(191,132)(181,132){1}
//: enddecls

  //: output g4 (Cout) @(274,142) /sn:0 /w:[ 0 ]
  and g8 (.I0(B), .I1(A), .Z(w13));   //: @(171,157) /sn:0 /delay:" 3" /w:[ 0 5 1 ]
  //: output g3 (S) @(272,100) /sn:0 /w:[ 0 ]
  //: input g2 (Cin) @(97,123) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(93,104) /sn:0 /w:[ 5 ]
  //: joint g10 (Cin) @(156, 123) /w:[ -1 2 1 4 ]
  xor g6 (.I0(w7), .I1(Cin), .Z(S));   //: @(181,98) /sn:0 /delay:" 4" /w:[ 3 3 1 ]
  and g7 (.I0(Cin), .I1(w7), .Z(w12));   //: @(171,132) /sn:0 /delay:" 3" /w:[ 5 0 1 ]
  or g9 (.I0(w12), .I1(w13), .Z(Cout));   //: @(223,142) /sn:0 /delay:" 3" /w:[ 0 0 1 ]
  //: joint g12 (A) @(104, 85) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(A), .I1(B), .Z(w7));   //: @(134,89) /sn:0 /delay:" 4" /w:[ 3 3 5 ]
  //: joint g11 (w7) @(149, 89) /w:[ 2 -1 4 1 ]
  //: input g0 (A) @(95,85) /sn:0 /w:[ 0 ]
  //: joint g13 (B) @(113, 104) /w:[ 1 2 4 -1 ]

endmodule

module main;    //: root_module
wire [15:0] w6;    //: /sn:0 {0}(403,573)(316,573)(316,571)(307,571){1}
wire w13;    //: /sn:0 {0}(491,620)(491,677)(476,677){1}
//: {2}(474,675)(474,667)(1187,667)(1187,312){3}
//: {4}(472,677)(-146,677)(-146,465){5}
//: {6}(-144,463)(-71,463)(-71,453)(-63,453){7}
//: {8}(-148,463)(-240,463){9}
wire [31:0] w16;    //: /sn:0 {0}(660,389)(708,389)(708,388)(756,388){1}
//: {2}(760,388)(830,388)(830,325)(866,325){3}
//: {4}(758,386)(758,376)(760,376)(760,304){5}
wire [4:0] w7;    //: /sn:0 {0}(250,515)(250,440)(280,440)(280,430){1}
//: {2}(282,428)(295,428){3}
//: {4}(278,428)(272,428)(272,387)(403,387){5}
wire w34;    //: /sn:0 {0}(590,284)(590,324)(539,324)(539,335){1}
wire [31:0] w4;    //: /sn:0 {0}(78,468)(84,468)(84,429)(101,429){1}
//: {2}(105,429)(183,429){3}
//: {4}(184,429)(207,429)(207,431)(231,431){5}
//: {6}(232,431)(242,431)(242,446)(190,446)(190,496)(146,496)(146,484)(143,484){7}
//: {8}(142,484)(131,484)(131,520)(249,520){9}
//: {10}(250,520)(259,520)(259,514)(295,514){11}
//: {12}(296,514)(331,514)(331,507)(343,507){13}
//: {14}(344,507)(354,507)(354,516)(343,516)(343,528)(321,528)(321,546)(303,546)(303,570){15}
//: {16}(303,571)(303,627){17}
//: {18}(103,431)(103,441)(101,441)(101,571){19}
wire w39;    //: /sn:0 {0}(428,0)(1323,0)(1323,254)(1378,254)(1378,242){1}
wire w25;    //: /sn:0 {0}(583,71)(583,99)(616,99){1}
wire [31:0] w3;    //: /sn:0 {0}(78,261)(130,261)(130,189)(545,189){1}
//: {2}(546,189)(652,189){3}
//: {4}(656,189)(827,189)(827,179){5}
//: {6}(829,177)(866,177){7}
//: {8}(827,175)(827,-32)(1106,-32){9}
//: {10}(654,187)(654,135)(683,135)(683,150){11}
wire [31:0] w22;    //: /sn:0 {0}(1053,176)(1096,176)(1096,83){1}
//: {2}(1098,81)(1117,81){3}
//: {4}(1096,79)(1096,-52)(1106,-52){5}
wire w36;    //: /sn:0 {0}(428,-39)(999,-39)(999,56)(1065,56){1}
wire w0;    //: /sn:0 {0}(428,-83)(564,-83)(564,226){1}
//: {2}(562,228)(500,228)(500,777){3}
//: {4}(564,230)(564,271)(567,271){5}
wire [5:0] w20;    //: /sn:0 {0}(199,64)(199,49)(184,49)(184,59){1}
//: {2}(186,61)(255,61){3}
//: {4}(184,63)(184,424){5}
wire [31:0] w30;    //: /sn:0 /dp:1 {0}(812,594)(812,559)(823,559)(823,544)(829,544){1}
wire [31:0] w29;    //: /sn:0 /dp:1 {0}(858,538)(863,538)(863,441){1}
//: {2}(865,439)(909,439)(909,441)(912,441){3}
//: {4}(861,439)(858,439)(858,358)(866,358){5}
wire w37;    //: /sn:0 {0}(428,-21)(1445,-21)(1445,324)(1226,324)(1226,312){1}
wire w42;    //: /sn:0 /dp:1 {0}(469,105)(469,123)(539,123)(539,106){1}
//: {2}(541,104)(580,104)(580,255){3}
//: {4}(539,102)(539,89)(428,89){5}
wire [5:0] w19;    //: /sn:0 {0}(546,184)(546,147)(627,147){1}
wire w18;    //: /sn:0 {0}(1086,59)(1122,59)(1122,-19){1}
wire w12;    //: /sn:0 /dp:1 {0}(453,335)(453,314)(647,314)(647,97)(637,97){1}
wire [31:0] w23;    //: /sn:0 {0}(1053,369)(1087,369){1}
//: {2}(1091,369)(1116,369)(1116,234){3}
//: {4}(1118,232)(1141,232)(1141,340)(1311,340)(1311,229)(1362,229){5}
//: {6}(1116,230)(1116,180)(1166,180){7}
//: {8}(1089,371)(1089,542)(1103,542)(1103,557)(1093,557){9}
wire [31:0] w10;    //: /sn:0 {0}(660,586)(666,586)(666,585)(673,585){1}
//: {2}(677,585)(717,585)(717,532){3}
//: {4}(719,530)(813,530)(813,532)(829,532){5}
//: {6}(717,528)(717,421)(737,421)(737,212)(866,212){7}
//: {8}(675,587)(675,810)(516,810){9}
wire w24;    //: /sn:0 {0}(1053,328)(1061,328)(1061,320){1}
//: {2}(1063,318)(1076,318)(1076,308){3}
//: {4}(1061,316)(1061,218){5}
//: {6}(1061,214)(1061,61)(1065,61){7}
//: {8}(1059,216)(600,216)(600,255){9}
wire w21;    //: /sn:0 {0}(603,71)(603,94)(616,94){1}
wire w1;    //: /sn:0 {0}(-63,303)(-110,303)(-110,688){1}
//: {2}(-108,690)(548,690)(548,620){3}
//: {4}(-112,690)(-232,690){5}
wire [31:0] w31;    //: /sn:0 /dp:1 {0}(424,620)(424,646)(473,646)(473,800)(487,800){1}
wire [31:0] w32;    //: /sn:0 {0}(1391,219)(1401,219)(1401,428){1}
//: {2}(1403,430)(1472,430)(1472,415){3}
//: {4}(1401,432)(1401,790)(516,790){5}
wire [4:0] w8;    //: /sn:0 {0}(403,487)(385,487)(385,486)(368,486){1}
//: {2}(364,486)(344,486)(344,502){3}
//: {4}(366,488)(366,498)(376,498)(376,723){5}
wire [31:0] w27;    //: /sn:0 /dp:1 {0}(633,152)(681,152)(681,-109)(1152,-109)(1152,-72)(1194,-72){1}
wire [3:0] w17;    //: /sn:0 {0}(428,23)(952,23)(952,85){1}
wire [31:0] w33;    //: /sn:0 {0}(1135,-42)(1184,-42)(1184,-52)(1194,-52){1}
wire [31:0] w28;    //: /sn:0 {0}(1296,164)(1354,164)(1354,180){1}
//: {2}(1356,182)(1565,182)(1565,129){3}
//: {4}(1354,184)(1354,209)(1362,209){5}
wire [31:0] w35;    //: /sn:0 {0}(1223,-62)(1239,-62)(1239,-157)(-73,-157)(-73,-24){1}
//: {2}(-75,-22)(-179,-22)(-179,-36){3}
//: {4}(-73,-20)(-73,380)(-63,380){5}
wire w14;    //: /sn:0 {0}(428,-57)(1081,-57)(1081,-134)(1179,-134)(1179,-27)(1210,-27)(1210,-39){1}
wire [31:0] w41;    //: /sn:0 {0}(893,614)(903,614)(903,599)(879,599)(879,571)(819,571)(819,556)(829,556){1}
wire [5:0] w2;    //: /sn:0 /dp:1 {0}(143,479)(143,-54)(255,-54){1}
wire w11;    //: /sn:0 {0}(428,-72)(456,-72)(456,309)(381,309)(381,516)(403,516){1}
wire [31:0] w15;    //: /sn:0 {0}(660,498)(704,498)(704,497)(749,497){1}
//: {2}(753,497)(811,497){3}
//: {4}(815,497)(1160,497)(1160,249)(1166,249){5}
//: {6}(813,499)(813,520)(829,520){7}
//: {8}(751,499)(751,509)(757,509)(757,727){9}
wire [25:0] w5;    //: /sn:0 /dp:1 {0}(627,157)(582,157)(582,129)(232,129)(232,426){1}
wire [4:0] w9;    //: /sn:0 /dp:1 {0}(296,509)(296,438)(403,438){1}
wire [1:0] w26;    //: /sn:0 /dp:5 {0}(845,561)(845,573)(774,573)(774,67)(603,67){1}
//: {2}(602,67)(583,67){3}
//: {4}(582,67)(428,67){5}
wire w40;    //: /sn:0 {0}(428,41)(1229,41)(1229,136){1}
//: enddecls

  concat g4 (.I0(w5), .I1(w19), .Z(w27));   //: @(632,152) /sn:0 /w:[ 0 1 0 ] /dr:0
  //: joint g44 (w20) @(184, 61) /w:[ 2 1 -1 4 ]
  tran g8(.Z(w9), .I(w4[20:16]));   //: @(296,512) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:0
  //: joint g3 (w28) @(1354, 182) /w:[ 2 1 -1 4 ]
  led g47 (.I(w22));   //: @(1124,81) /sn:0 /R:3 /w:[ 3 ] /type:2
  //: joint g16 (w15) @(813, 497) /w:[ 4 -1 3 6 ]
  //: joint g26 (w16) @(758, 388) /w:[ 2 4 1 -1 ]
  //: joint g17 (w3) @(827, 177) /w:[ 6 8 -1 5 ]
  EXE g2 (.ALU_operation(w17), .data_read_2(w29), .data_read_1(w16), .PCNext(w3), .INM32(w10), .Zero_signal(w24), .ALU_result(w23), .branch_target(w22));   //: @(867, 86) /sz:(185, 314) /sn:0 /p:[ Ti0>1 Li0>5 Li1>3 Li2>7 Li3>7 Ro0<0 Ro1<0 Ro2<0 ]
  led g30 (.I(w35));   //: @(-179,-43) /sn:0 /w:[ 3 ] /type:2
  and g23 (.I0(w36), .I1(w24), .Z(w18));   //: @(1076,59) /sn:0 /w:[ 1 7 0 ]
  led g24 (.I(w16));   //: @(760,297) /sn:0 /w:[ 5 ] /type:2
  //: joint g39 (w15) @(751, 497) /w:[ 2 -1 1 8 ]
  READ g1 (.Pop(w12), .RegWrite(w34), .Read_register_1(w7), .Read_register_2(w9), .Write_register(w8), .mux_RegDst(w11), .Sign_ext_in(w6), .clk(w13), .clr(w1), .Write_data(w31), .Read_data_1(w16), .Read_data_2(w15), .Sign_ext_out(w10));   //: @(404, 336) /sz:(255, 283) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>5 Li1>1 Li2>0 Li3>1 Li4>0 Bi0>0 Bi1>3 Bi2>0 Ro0<0 Ro1<0 Ro2<0 ]
  //: joint g29 (w4) @(103, 429) /w:[ 2 -1 1 18 ]
  tran g60(.Z(w25), .I(w26[1]));   //: @(583,65) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  led g51 (.I(w24));   //: @(1076,301) /sn:0 /w:[ 3 ] /type:0
  ctrl ctrl (.funct(w20), .op(w2), .cmpseti(w0), .RegWrite(w42), .ALUSrc(w26), .MemWrite(w40), .MemtoReg(w39), .ALUCtrl(w17), .MemRead(w37), .Branch(w36), .Jump(w14), .RegDst(w11));   //: @(256, -88) /sz:(171, 204) /sn:0 /p:[ Li0>3 Li1>1 Ro0<0 Ro1<5 Ro2<5 Ro3<0 Ro4<0 Ro5<0 Ro6<0 Ro7<0 Ro8<0 Ro9<0 ]
  mux g18 (.I0(w33), .I1(w27), .S(w14), .Z(w35));   //: @(1210,-62) /sn:0 /R:1 /w:[ 1 1 1 0 ] /ss:0 /do:0
  tran g10(.Z(w6), .I(w4[15:0]));   //: @(301,571) /sn:0 /R:2 /w:[ 1 16 15 ] /ss:1
  //: joint g25 (w13) @(-146, 463) /w:[ 6 -1 8 5 ]
  mux g49 (.I0(w42), .I1(w24), .S(w0), .Z(w34));   //: @(590,271) /sn:0 /w:[ 3 9 5 0 ] /ss:0 /do:0
  tran g6(.Z(w5), .I(w4[25:0]));   //: @(232,429) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:0
  //: joint g50 (w42) @(539, 104) /w:[ 2 4 -1 1 ]
  //: joint g35 (w23) @(1089, 369) /w:[ 2 -1 1 8 ]
  tran g7(.Z(w7), .I(w4[25:21]));   //: @(250,518) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:0
  tran g9(.Z(w8), .I(w4[15:11]));   //: @(344,505) /sn:0 /R:1 /w:[ 3 13 14 ] /ss:0
  //: joint g56 (w0) @(564, 228) /w:[ -1 1 2 4 ]
  tran g58(.Z(w21), .I(w26[0]));   //: @(603,65) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  led g59 (.I(w42));   //: @(469,98) /sn:0 /w:[ 0 ] /type:0
  MEM Mem (.memWrite(w40), .Address(w23), .write_data(w15), .clk(w13), .MemRead(w37), .read_data(w28));   //: @(1167, 137) /sz:(128, 174) /sn:0 /p:[ Ti0>1 Li0>7 Li1>5 Bi0>3 Bi1>1 Ro0<0 ]
  //: joint g31 (w35) @(-73, -22) /w:[ -1 1 2 4 ]
  tran g22(.Z(w2), .I(w4[31:26]));   //: @(143,482) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:0
  //: joint g54 (w8) @(366, 486) /w:[ 1 -1 2 4 ]
  led g36 (.I(w3));   //: @(683,157) /sn:0 /R:2 /w:[ 11 ] /type:2
  //: joint g45 (w29) @(863, 439) /w:[ 2 -1 4 1 ]
  mux g41 (.I0(w32), .I1(w10), .S(w0), .Z(w31));   //: @(500,800) /sn:0 /R:3 /w:[ 5 9 3 1 ] /ss:0 /do:0
  //: joint g33 (w10) @(675, 585) /w:[ 2 -1 1 8 ]
  //: joint g52 (w24) @(1061, 318) /w:[ 2 4 -1 1 ]
  //: joint g40 (w13) @(474, 677) /w:[ 1 2 4 -1 ]
  //: dip g42 (w30) @(812,605) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: joint g12 (w10) @(717, 530) /w:[ 4 6 -1 3 ]
  clock clk (.Z(w13));   //: @(-253,463) /sn:0 /w:[ 9 ] /omega:2000 /phi:0 /duty:50
  led g34 (.I(w23));   //: @(1086,557) /sn:0 /R:1 /w:[ 9 ] /type:2
  led g28 (.I(w4));   //: @(101,578) /sn:0 /R:2 /w:[ 19 ] /type:2
  //: joint g46 (w32) @(1401, 430) /w:[ 2 1 -1 4 ]
  and g57 (.I0(w21), .I1(w25), .Z(w12));   //: @(627,97) /sn:0 /w:[ 1 1 1 ]
  //: switch g11 (w41) @(876,614) /sn:0 /w:[ 0 ] /st:0
  tran g5(.Z(w19), .I(w3[31:26]));   //: @(546,187) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0
  //: joint g14 (w23) @(1116, 232) /w:[ 4 6 -1 3 ]
  //: joint g19 (w7) @(280, 428) /w:[ 2 -1 4 1 ]
  tran g21(.Z(w20), .I(w4[5:0]));   //: @(184,427) /sn:0 /R:1 /w:[ 5 3 4 ] /ss:0
  //: switch reset (w1) @(-249,690) /sn:0 /w:[ 5 ] /st:0
  fetch Fetch (.PCNew(w35), .reset(w1), .clk(w13), .Inst(w4), .PCNext(w3));   //: @(-62, 217) /sz:(139, 319) /sn:0 /p:[ Li0>5 Li1>0 Li2>7 Ro0<0 Ro1<0 ]
  led g32 (.I(w32));   //: @(1472,408) /sn:0 /w:[ 3 ] /type:2
  mux g20 (.I0(w15), .I1(w10), .I2(w30), .I3(w41), .S(w26), .Z(w29));   //: @(845,538) /sn:0 /R:1 /w:[ 7 5 1 1 0 0 ] /ss:0 /do:1
  led g0 (.I(w28));   //: @(1565,122) /sn:0 /w:[ 3 ] /type:2
  led g38 (.I(w15));   //: @(757,734) /sn:0 /R:2 /w:[ 9 ] /type:2
  mux g15 (.I0(w3), .I1(w22), .S(w18), .Z(w33));   //: @(1122,-42) /sn:0 /R:1 /w:[ 9 5 1 0 ] /ss:0 /do:0
  led g43 (.I(w29));   //: @(919,441) /sn:0 /R:3 /w:[ 3 ] /type:2
  //: joint g27 (w1) @(-110, 690) /w:[ 2 1 4 -1 ]
  //: joint g48 (w22) @(1096, 81) /w:[ 2 4 -1 1 ]
  //: joint g37 (w3) @(654, 189) /w:[ 4 10 3 -1 ]
  //: joint g55 (w24) @(1061, 216) /w:[ -1 6 8 5 ]
  led g53 (.I(w8));   //: @(376,730) /sn:0 /R:2 /w:[ 5 ] /type:2
  mux g13 (.I0(w23), .I1(w28), .S(w39), .Z(w32));   //: @(1378,219) /sn:0 /R:1 /w:[ 5 5 1 0 ] /ss:0 /do:0

endmodule

module CLA(A, S, B, Cin, g0, p0);
//: interface  /sz:(162, 96) /bd:[ Ti0>B[3:0](61/162) Ti1>A[3:0](24/162) Ti2>B[3:0](61/162) Ti3>A[3:0](24/162) Ri0>Cin(34/96) Ri1>Cin(34/96) Bo0<p0(130/162) Bo1<g0(87/162) Bo2<S[3:0](24/162) Bo3<p0(130/162) Bo4<g0(87/162) Bo5<S[3:0](24/162) ]
input [3:0] B;    //: /sn:0 {0}(117,75)(205,75){1}
//: {2}(206,75)(306,75){3}
//: {4}(307,75)(406,75){5}
//: {6}(407,75)(498,75){7}
//: {8}(499,75)(559,75){9}
input [3:0] A;    //: /sn:0 {0}(126,58)(175,58){1}
//: {2}(176,58)(277,58){3}
//: {4}(278,58)(378,58){5}
//: {6}(379,58)(469,58){7}
//: {8}(470,58)(557,58){9}
input Cin;    //: /sn:0 {0}(574,109)(557,109){1}
//: {2}(553,109)(526,109)(526,120){3}
//: {4}(555,111)(555,238)(538,238){5}
output p0;    //: /sn:0 {0}(483,306)(493,306)(493,292)(474,292)(474,267)(483,267)(483,257){1}
output g0;    //: /sn:0 {0}(432,303)(422,303)(422,288)(458,288)(458,257){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(639,197)(721,197){1}
wire w6;    //: /sn:0 {0}(278,123)(278,62){1}
wire w13;    //: /sn:0 {0}(407,122)(407,79){1}
wire w16;    //: /sn:0 {0}(412,164)(412,205)(413,205)(413,215){1}
wire w7;    //: /sn:0 {0}(307,123)(307,79){1}
wire w4;    //: /sn:0 {0}(201,164)(201,215){1}
wire w0;    //: /sn:0 {0}(176,122)(176,62){1}
wire w3;    //: /sn:0 {0}(174,164)(174,182)(633,182){1}
wire w22;    //: /sn:0 {0}(505,165)(505,205)(504,205)(504,215){1}
wire w20;    //: /sn:0 /dp:1 {0}(448,215)(448,112)(433,112)(433,122){1}
wire w12;    //: /sn:0 {0}(379,122)(379,62){1}
wire w18;    //: /sn:0 {0}(470,120)(470,62){1}
wire w19;    //: /sn:0 {0}(499,120)(499,79){1}
wire w10;    //: /sn:0 {0}(313,165)(313,215){1}
wire w23;    //: /sn:0 {0}(526,165)(526,205)(527,205)(527,215){1}
wire w21;    //: /sn:0 {0}(478,165)(478,212)(633,212){1}
wire w1;    //: /sn:0 {0}(206,122)(206,79){1}
wire w8;    //: /sn:0 /dp:1 {0}(250,215)(250,112)(234,112)(234,122){1}
wire w17;    //: /sn:0 {0}(433,164)(433,205)(434,205)(434,215){1}
wire w14;    //: /sn:0 /dp:1 {0}(353,215)(353,113)(334,113)(334,123){1}
wire w11;    //: /sn:0 {0}(334,165)(334,205)(335,205)(335,215){1}
wire w2;    //: /sn:0 {0}(143,237)(153,237){1}
wire w15;    //: /sn:0 {0}(386,164)(386,202)(633,202){1}
wire w5;    //: /sn:0 {0}(225,164)(225,205)(226,205)(226,215){1}
wire w9;    //: /sn:0 {0}(286,165)(286,192)(633,192){1}
//: enddecls

  //: input g4 (A) @(559,58) /sn:0 /R:2 /w:[ 9 ]
  tran g8(.Z(w0), .I(A[3]));   //: @(176,56) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  PFA g3 (.Ci(Cin), .B(w19), .A(w18), .Gi(w23), .Pi(w22), .S(w21));   //: @(455, 121) /sz:(77, 43) /sn:0 /p:[ Ti0>3 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  CLL g16 (.P3(w4), .G3(w5), .P2(w10), .G2(w11), .P1(w16), .G1(w17), .P0(w22), .G0(w23), .Cin(Cin), .C3(w8), .C2(w14), .C1(w20), .C4(w2), .PG(p0), .GG(g0));   //: @(154, 216) /sz:(383, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>5 To0<0 To1<0 To2<0 Lo0<1 Bo0<1 Bo1<1 ]
  concat g17 (.I0(w21), .I1(w15), .I2(w9), .I3(w3), .Z(S));   //: @(638,197) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  PFA g2 (.Ci(w20), .B(w13), .A(w12), .Gi(w17), .Pi(w16), .S(w15));   //: @(364, 123) /sz:(75, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  PFA g1 (.Ci(w14), .B(w7), .A(w6), .Gi(w11), .Pi(w10), .S(w9));   //: @(263, 124) /sz:(77, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  //: output g18 (S) @(718,197) /sn:0 /w:[ 1 ]
  tran g10(.Z(w19), .I(B[0]));   //: @(499,73) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g6(.Z(w12), .I(A[1]));   //: @(379,56) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g7(.Z(w6), .I(A[2]));   //: @(278,56) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: input g9 (B) @(561,75) /sn:0 /R:2 /w:[ 9 ]
  tran g12(.Z(w7), .I(B[2]));   //: @(307,73) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g5(.Z(w18), .I(A[0]));   //: @(470,56) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g11(.Z(w13), .I(B[1]));   //: @(407,73) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g14 (Cin) @(576,109) /sn:0 /R:2 /w:[ 0 ]
  //: output g19 (g0) @(429,303) /sn:0 /w:[ 0 ]
  //: output g20 (p0) @(486,306) /sn:0 /R:2 /w:[ 0 ]
  PFA g0 (.Ci(w8), .B(w1), .A(w0), .Gi(w5), .Pi(w4), .S(w3));   //: @(160, 123) /sz:(80, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  //: joint g15 (Cin) @(555, 109) /w:[ 1 -1 2 4 ]
  tran g13(.Z(w1), .I(B[3]));   //: @(206,73) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1

endmodule
